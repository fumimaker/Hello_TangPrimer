// Verilog netlist created by TD v4.6.14756
// Thu Mar 12 20:59:10 2020

`timescale 1ns / 1ps
module bitmaprom  // al_ip/bitmaprom.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [15:0] addra;  // al_ip/bitmaprom.v(18)
  input clka;  // al_ip/bitmaprom.v(19)
  input rsta;  // al_ip/bitmaprom.v(20)
  output [8:0] doa;  // al_ip/bitmaprom.v(16)

  wire [0:5] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b0/B0_10 ;
  wire  \inst_doa_mux_b0/B0_11 ;
  wire  \inst_doa_mux_b0/B0_12 ;
  wire  \inst_doa_mux_b0/B0_13 ;
  wire  \inst_doa_mux_b0/B0_14 ;
  wire  \inst_doa_mux_b0/B0_15 ;
  wire  \inst_doa_mux_b0/B0_16 ;
  wire  \inst_doa_mux_b0/B0_17 ;
  wire  \inst_doa_mux_b0/B0_18 ;
  wire  \inst_doa_mux_b0/B0_19 ;
  wire  \inst_doa_mux_b0/B0_2 ;
  wire  \inst_doa_mux_b0/B0_20 ;
  wire  \inst_doa_mux_b0/B0_21 ;
  wire  \inst_doa_mux_b0/B0_22 ;
  wire  \inst_doa_mux_b0/B0_23 ;
  wire  \inst_doa_mux_b0/B0_24 ;
  wire  \inst_doa_mux_b0/B0_25 ;
  wire  \inst_doa_mux_b0/B0_26 ;
  wire  \inst_doa_mux_b0/B0_27 ;
  wire  \inst_doa_mux_b0/B0_28 ;
  wire  \inst_doa_mux_b0/B0_29 ;
  wire  \inst_doa_mux_b0/B0_3 ;
  wire  \inst_doa_mux_b0/B0_30 ;
  wire  \inst_doa_mux_b0/B0_31 ;
  wire  \inst_doa_mux_b0/B0_4 ;
  wire  \inst_doa_mux_b0/B0_5 ;
  wire  \inst_doa_mux_b0/B0_6 ;
  wire  \inst_doa_mux_b0/B0_7 ;
  wire  \inst_doa_mux_b0/B0_8 ;
  wire  \inst_doa_mux_b0/B0_9 ;
  wire  \inst_doa_mux_b0/B1_0 ;
  wire  \inst_doa_mux_b0/B1_1 ;
  wire  \inst_doa_mux_b0/B1_10 ;
  wire  \inst_doa_mux_b0/B1_11 ;
  wire  \inst_doa_mux_b0/B1_12 ;
  wire  \inst_doa_mux_b0/B1_13 ;
  wire  \inst_doa_mux_b0/B1_14 ;
  wire  \inst_doa_mux_b0/B1_15 ;
  wire  \inst_doa_mux_b0/B1_2 ;
  wire  \inst_doa_mux_b0/B1_3 ;
  wire  \inst_doa_mux_b0/B1_4 ;
  wire  \inst_doa_mux_b0/B1_5 ;
  wire  \inst_doa_mux_b0/B1_6 ;
  wire  \inst_doa_mux_b0/B1_7 ;
  wire  \inst_doa_mux_b0/B1_8 ;
  wire  \inst_doa_mux_b0/B1_9 ;
  wire  \inst_doa_mux_b0/B2_0 ;
  wire  \inst_doa_mux_b0/B2_1 ;
  wire  \inst_doa_mux_b0/B2_2 ;
  wire  \inst_doa_mux_b0/B2_3 ;
  wire  \inst_doa_mux_b0/B2_4 ;
  wire  \inst_doa_mux_b0/B2_5 ;
  wire  \inst_doa_mux_b0/B2_6 ;
  wire  \inst_doa_mux_b0/B2_7 ;
  wire  \inst_doa_mux_b0/B3_0 ;
  wire  \inst_doa_mux_b0/B3_1 ;
  wire  \inst_doa_mux_b0/B3_2 ;
  wire  \inst_doa_mux_b0/B3_3 ;
  wire  \inst_doa_mux_b0/B4_0 ;
  wire  \inst_doa_mux_b0/B4_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b1/B0_10 ;
  wire  \inst_doa_mux_b1/B0_11 ;
  wire  \inst_doa_mux_b1/B0_12 ;
  wire  \inst_doa_mux_b1/B0_13 ;
  wire  \inst_doa_mux_b1/B0_14 ;
  wire  \inst_doa_mux_b1/B0_15 ;
  wire  \inst_doa_mux_b1/B0_16 ;
  wire  \inst_doa_mux_b1/B0_17 ;
  wire  \inst_doa_mux_b1/B0_18 ;
  wire  \inst_doa_mux_b1/B0_19 ;
  wire  \inst_doa_mux_b1/B0_2 ;
  wire  \inst_doa_mux_b1/B0_20 ;
  wire  \inst_doa_mux_b1/B0_21 ;
  wire  \inst_doa_mux_b1/B0_22 ;
  wire  \inst_doa_mux_b1/B0_23 ;
  wire  \inst_doa_mux_b1/B0_24 ;
  wire  \inst_doa_mux_b1/B0_25 ;
  wire  \inst_doa_mux_b1/B0_26 ;
  wire  \inst_doa_mux_b1/B0_27 ;
  wire  \inst_doa_mux_b1/B0_28 ;
  wire  \inst_doa_mux_b1/B0_29 ;
  wire  \inst_doa_mux_b1/B0_3 ;
  wire  \inst_doa_mux_b1/B0_30 ;
  wire  \inst_doa_mux_b1/B0_31 ;
  wire  \inst_doa_mux_b1/B0_4 ;
  wire  \inst_doa_mux_b1/B0_5 ;
  wire  \inst_doa_mux_b1/B0_6 ;
  wire  \inst_doa_mux_b1/B0_7 ;
  wire  \inst_doa_mux_b1/B0_8 ;
  wire  \inst_doa_mux_b1/B0_9 ;
  wire  \inst_doa_mux_b1/B1_0 ;
  wire  \inst_doa_mux_b1/B1_1 ;
  wire  \inst_doa_mux_b1/B1_10 ;
  wire  \inst_doa_mux_b1/B1_11 ;
  wire  \inst_doa_mux_b1/B1_12 ;
  wire  \inst_doa_mux_b1/B1_13 ;
  wire  \inst_doa_mux_b1/B1_14 ;
  wire  \inst_doa_mux_b1/B1_15 ;
  wire  \inst_doa_mux_b1/B1_2 ;
  wire  \inst_doa_mux_b1/B1_3 ;
  wire  \inst_doa_mux_b1/B1_4 ;
  wire  \inst_doa_mux_b1/B1_5 ;
  wire  \inst_doa_mux_b1/B1_6 ;
  wire  \inst_doa_mux_b1/B1_7 ;
  wire  \inst_doa_mux_b1/B1_8 ;
  wire  \inst_doa_mux_b1/B1_9 ;
  wire  \inst_doa_mux_b1/B2_0 ;
  wire  \inst_doa_mux_b1/B2_1 ;
  wire  \inst_doa_mux_b1/B2_2 ;
  wire  \inst_doa_mux_b1/B2_3 ;
  wire  \inst_doa_mux_b1/B2_4 ;
  wire  \inst_doa_mux_b1/B2_5 ;
  wire  \inst_doa_mux_b1/B2_6 ;
  wire  \inst_doa_mux_b1/B2_7 ;
  wire  \inst_doa_mux_b1/B3_0 ;
  wire  \inst_doa_mux_b1/B3_1 ;
  wire  \inst_doa_mux_b1/B3_2 ;
  wire  \inst_doa_mux_b1/B3_3 ;
  wire  \inst_doa_mux_b1/B4_0 ;
  wire  \inst_doa_mux_b1/B4_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b2/B0_10 ;
  wire  \inst_doa_mux_b2/B0_11 ;
  wire  \inst_doa_mux_b2/B0_12 ;
  wire  \inst_doa_mux_b2/B0_13 ;
  wire  \inst_doa_mux_b2/B0_14 ;
  wire  \inst_doa_mux_b2/B0_15 ;
  wire  \inst_doa_mux_b2/B0_16 ;
  wire  \inst_doa_mux_b2/B0_17 ;
  wire  \inst_doa_mux_b2/B0_18 ;
  wire  \inst_doa_mux_b2/B0_19 ;
  wire  \inst_doa_mux_b2/B0_2 ;
  wire  \inst_doa_mux_b2/B0_20 ;
  wire  \inst_doa_mux_b2/B0_21 ;
  wire  \inst_doa_mux_b2/B0_22 ;
  wire  \inst_doa_mux_b2/B0_23 ;
  wire  \inst_doa_mux_b2/B0_24 ;
  wire  \inst_doa_mux_b2/B0_25 ;
  wire  \inst_doa_mux_b2/B0_26 ;
  wire  \inst_doa_mux_b2/B0_27 ;
  wire  \inst_doa_mux_b2/B0_28 ;
  wire  \inst_doa_mux_b2/B0_29 ;
  wire  \inst_doa_mux_b2/B0_3 ;
  wire  \inst_doa_mux_b2/B0_30 ;
  wire  \inst_doa_mux_b2/B0_31 ;
  wire  \inst_doa_mux_b2/B0_4 ;
  wire  \inst_doa_mux_b2/B0_5 ;
  wire  \inst_doa_mux_b2/B0_6 ;
  wire  \inst_doa_mux_b2/B0_7 ;
  wire  \inst_doa_mux_b2/B0_8 ;
  wire  \inst_doa_mux_b2/B0_9 ;
  wire  \inst_doa_mux_b2/B1_0 ;
  wire  \inst_doa_mux_b2/B1_1 ;
  wire  \inst_doa_mux_b2/B1_10 ;
  wire  \inst_doa_mux_b2/B1_11 ;
  wire  \inst_doa_mux_b2/B1_12 ;
  wire  \inst_doa_mux_b2/B1_13 ;
  wire  \inst_doa_mux_b2/B1_14 ;
  wire  \inst_doa_mux_b2/B1_15 ;
  wire  \inst_doa_mux_b2/B1_2 ;
  wire  \inst_doa_mux_b2/B1_3 ;
  wire  \inst_doa_mux_b2/B1_4 ;
  wire  \inst_doa_mux_b2/B1_5 ;
  wire  \inst_doa_mux_b2/B1_6 ;
  wire  \inst_doa_mux_b2/B1_7 ;
  wire  \inst_doa_mux_b2/B1_8 ;
  wire  \inst_doa_mux_b2/B1_9 ;
  wire  \inst_doa_mux_b2/B2_0 ;
  wire  \inst_doa_mux_b2/B2_1 ;
  wire  \inst_doa_mux_b2/B2_2 ;
  wire  \inst_doa_mux_b2/B2_3 ;
  wire  \inst_doa_mux_b2/B2_4 ;
  wire  \inst_doa_mux_b2/B2_5 ;
  wire  \inst_doa_mux_b2/B2_6 ;
  wire  \inst_doa_mux_b2/B2_7 ;
  wire  \inst_doa_mux_b2/B3_0 ;
  wire  \inst_doa_mux_b2/B3_1 ;
  wire  \inst_doa_mux_b2/B3_2 ;
  wire  \inst_doa_mux_b2/B3_3 ;
  wire  \inst_doa_mux_b2/B4_0 ;
  wire  \inst_doa_mux_b2/B4_1 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b3/B0_10 ;
  wire  \inst_doa_mux_b3/B0_11 ;
  wire  \inst_doa_mux_b3/B0_12 ;
  wire  \inst_doa_mux_b3/B0_13 ;
  wire  \inst_doa_mux_b3/B0_14 ;
  wire  \inst_doa_mux_b3/B0_15 ;
  wire  \inst_doa_mux_b3/B0_16 ;
  wire  \inst_doa_mux_b3/B0_17 ;
  wire  \inst_doa_mux_b3/B0_18 ;
  wire  \inst_doa_mux_b3/B0_19 ;
  wire  \inst_doa_mux_b3/B0_2 ;
  wire  \inst_doa_mux_b3/B0_20 ;
  wire  \inst_doa_mux_b3/B0_21 ;
  wire  \inst_doa_mux_b3/B0_22 ;
  wire  \inst_doa_mux_b3/B0_23 ;
  wire  \inst_doa_mux_b3/B0_24 ;
  wire  \inst_doa_mux_b3/B0_25 ;
  wire  \inst_doa_mux_b3/B0_26 ;
  wire  \inst_doa_mux_b3/B0_27 ;
  wire  \inst_doa_mux_b3/B0_28 ;
  wire  \inst_doa_mux_b3/B0_29 ;
  wire  \inst_doa_mux_b3/B0_3 ;
  wire  \inst_doa_mux_b3/B0_30 ;
  wire  \inst_doa_mux_b3/B0_31 ;
  wire  \inst_doa_mux_b3/B0_4 ;
  wire  \inst_doa_mux_b3/B0_5 ;
  wire  \inst_doa_mux_b3/B0_6 ;
  wire  \inst_doa_mux_b3/B0_7 ;
  wire  \inst_doa_mux_b3/B0_8 ;
  wire  \inst_doa_mux_b3/B0_9 ;
  wire  \inst_doa_mux_b3/B1_0 ;
  wire  \inst_doa_mux_b3/B1_1 ;
  wire  \inst_doa_mux_b3/B1_10 ;
  wire  \inst_doa_mux_b3/B1_11 ;
  wire  \inst_doa_mux_b3/B1_12 ;
  wire  \inst_doa_mux_b3/B1_13 ;
  wire  \inst_doa_mux_b3/B1_14 ;
  wire  \inst_doa_mux_b3/B1_15 ;
  wire  \inst_doa_mux_b3/B1_2 ;
  wire  \inst_doa_mux_b3/B1_3 ;
  wire  \inst_doa_mux_b3/B1_4 ;
  wire  \inst_doa_mux_b3/B1_5 ;
  wire  \inst_doa_mux_b3/B1_6 ;
  wire  \inst_doa_mux_b3/B1_7 ;
  wire  \inst_doa_mux_b3/B1_8 ;
  wire  \inst_doa_mux_b3/B1_9 ;
  wire  \inst_doa_mux_b3/B2_0 ;
  wire  \inst_doa_mux_b3/B2_1 ;
  wire  \inst_doa_mux_b3/B2_2 ;
  wire  \inst_doa_mux_b3/B2_3 ;
  wire  \inst_doa_mux_b3/B2_4 ;
  wire  \inst_doa_mux_b3/B2_5 ;
  wire  \inst_doa_mux_b3/B2_6 ;
  wire  \inst_doa_mux_b3/B2_7 ;
  wire  \inst_doa_mux_b3/B3_0 ;
  wire  \inst_doa_mux_b3/B3_1 ;
  wire  \inst_doa_mux_b3/B3_2 ;
  wire  \inst_doa_mux_b3/B3_3 ;
  wire  \inst_doa_mux_b3/B4_0 ;
  wire  \inst_doa_mux_b3/B4_1 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b4/B0_10 ;
  wire  \inst_doa_mux_b4/B0_11 ;
  wire  \inst_doa_mux_b4/B0_12 ;
  wire  \inst_doa_mux_b4/B0_13 ;
  wire  \inst_doa_mux_b4/B0_14 ;
  wire  \inst_doa_mux_b4/B0_15 ;
  wire  \inst_doa_mux_b4/B0_16 ;
  wire  \inst_doa_mux_b4/B0_17 ;
  wire  \inst_doa_mux_b4/B0_18 ;
  wire  \inst_doa_mux_b4/B0_19 ;
  wire  \inst_doa_mux_b4/B0_2 ;
  wire  \inst_doa_mux_b4/B0_20 ;
  wire  \inst_doa_mux_b4/B0_21 ;
  wire  \inst_doa_mux_b4/B0_22 ;
  wire  \inst_doa_mux_b4/B0_23 ;
  wire  \inst_doa_mux_b4/B0_24 ;
  wire  \inst_doa_mux_b4/B0_25 ;
  wire  \inst_doa_mux_b4/B0_26 ;
  wire  \inst_doa_mux_b4/B0_27 ;
  wire  \inst_doa_mux_b4/B0_28 ;
  wire  \inst_doa_mux_b4/B0_29 ;
  wire  \inst_doa_mux_b4/B0_3 ;
  wire  \inst_doa_mux_b4/B0_30 ;
  wire  \inst_doa_mux_b4/B0_31 ;
  wire  \inst_doa_mux_b4/B0_4 ;
  wire  \inst_doa_mux_b4/B0_5 ;
  wire  \inst_doa_mux_b4/B0_6 ;
  wire  \inst_doa_mux_b4/B0_7 ;
  wire  \inst_doa_mux_b4/B0_8 ;
  wire  \inst_doa_mux_b4/B0_9 ;
  wire  \inst_doa_mux_b4/B1_0 ;
  wire  \inst_doa_mux_b4/B1_1 ;
  wire  \inst_doa_mux_b4/B1_10 ;
  wire  \inst_doa_mux_b4/B1_11 ;
  wire  \inst_doa_mux_b4/B1_12 ;
  wire  \inst_doa_mux_b4/B1_13 ;
  wire  \inst_doa_mux_b4/B1_14 ;
  wire  \inst_doa_mux_b4/B1_15 ;
  wire  \inst_doa_mux_b4/B1_2 ;
  wire  \inst_doa_mux_b4/B1_3 ;
  wire  \inst_doa_mux_b4/B1_4 ;
  wire  \inst_doa_mux_b4/B1_5 ;
  wire  \inst_doa_mux_b4/B1_6 ;
  wire  \inst_doa_mux_b4/B1_7 ;
  wire  \inst_doa_mux_b4/B1_8 ;
  wire  \inst_doa_mux_b4/B1_9 ;
  wire  \inst_doa_mux_b4/B2_0 ;
  wire  \inst_doa_mux_b4/B2_1 ;
  wire  \inst_doa_mux_b4/B2_2 ;
  wire  \inst_doa_mux_b4/B2_3 ;
  wire  \inst_doa_mux_b4/B2_4 ;
  wire  \inst_doa_mux_b4/B2_5 ;
  wire  \inst_doa_mux_b4/B2_6 ;
  wire  \inst_doa_mux_b4/B2_7 ;
  wire  \inst_doa_mux_b4/B3_0 ;
  wire  \inst_doa_mux_b4/B3_1 ;
  wire  \inst_doa_mux_b4/B3_2 ;
  wire  \inst_doa_mux_b4/B3_3 ;
  wire  \inst_doa_mux_b4/B4_0 ;
  wire  \inst_doa_mux_b4/B4_1 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b5/B0_10 ;
  wire  \inst_doa_mux_b5/B0_11 ;
  wire  \inst_doa_mux_b5/B0_12 ;
  wire  \inst_doa_mux_b5/B0_13 ;
  wire  \inst_doa_mux_b5/B0_14 ;
  wire  \inst_doa_mux_b5/B0_15 ;
  wire  \inst_doa_mux_b5/B0_16 ;
  wire  \inst_doa_mux_b5/B0_17 ;
  wire  \inst_doa_mux_b5/B0_18 ;
  wire  \inst_doa_mux_b5/B0_19 ;
  wire  \inst_doa_mux_b5/B0_2 ;
  wire  \inst_doa_mux_b5/B0_20 ;
  wire  \inst_doa_mux_b5/B0_21 ;
  wire  \inst_doa_mux_b5/B0_22 ;
  wire  \inst_doa_mux_b5/B0_23 ;
  wire  \inst_doa_mux_b5/B0_24 ;
  wire  \inst_doa_mux_b5/B0_25 ;
  wire  \inst_doa_mux_b5/B0_26 ;
  wire  \inst_doa_mux_b5/B0_27 ;
  wire  \inst_doa_mux_b5/B0_28 ;
  wire  \inst_doa_mux_b5/B0_29 ;
  wire  \inst_doa_mux_b5/B0_3 ;
  wire  \inst_doa_mux_b5/B0_30 ;
  wire  \inst_doa_mux_b5/B0_31 ;
  wire  \inst_doa_mux_b5/B0_4 ;
  wire  \inst_doa_mux_b5/B0_5 ;
  wire  \inst_doa_mux_b5/B0_6 ;
  wire  \inst_doa_mux_b5/B0_7 ;
  wire  \inst_doa_mux_b5/B0_8 ;
  wire  \inst_doa_mux_b5/B0_9 ;
  wire  \inst_doa_mux_b5/B1_0 ;
  wire  \inst_doa_mux_b5/B1_1 ;
  wire  \inst_doa_mux_b5/B1_10 ;
  wire  \inst_doa_mux_b5/B1_11 ;
  wire  \inst_doa_mux_b5/B1_12 ;
  wire  \inst_doa_mux_b5/B1_13 ;
  wire  \inst_doa_mux_b5/B1_14 ;
  wire  \inst_doa_mux_b5/B1_15 ;
  wire  \inst_doa_mux_b5/B1_2 ;
  wire  \inst_doa_mux_b5/B1_3 ;
  wire  \inst_doa_mux_b5/B1_4 ;
  wire  \inst_doa_mux_b5/B1_5 ;
  wire  \inst_doa_mux_b5/B1_6 ;
  wire  \inst_doa_mux_b5/B1_7 ;
  wire  \inst_doa_mux_b5/B1_8 ;
  wire  \inst_doa_mux_b5/B1_9 ;
  wire  \inst_doa_mux_b5/B2_0 ;
  wire  \inst_doa_mux_b5/B2_1 ;
  wire  \inst_doa_mux_b5/B2_2 ;
  wire  \inst_doa_mux_b5/B2_3 ;
  wire  \inst_doa_mux_b5/B2_4 ;
  wire  \inst_doa_mux_b5/B2_5 ;
  wire  \inst_doa_mux_b5/B2_6 ;
  wire  \inst_doa_mux_b5/B2_7 ;
  wire  \inst_doa_mux_b5/B3_0 ;
  wire  \inst_doa_mux_b5/B3_1 ;
  wire  \inst_doa_mux_b5/B3_2 ;
  wire  \inst_doa_mux_b5/B3_3 ;
  wire  \inst_doa_mux_b5/B4_0 ;
  wire  \inst_doa_mux_b5/B4_1 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b6/B0_10 ;
  wire  \inst_doa_mux_b6/B0_11 ;
  wire  \inst_doa_mux_b6/B0_12 ;
  wire  \inst_doa_mux_b6/B0_13 ;
  wire  \inst_doa_mux_b6/B0_14 ;
  wire  \inst_doa_mux_b6/B0_15 ;
  wire  \inst_doa_mux_b6/B0_16 ;
  wire  \inst_doa_mux_b6/B0_17 ;
  wire  \inst_doa_mux_b6/B0_18 ;
  wire  \inst_doa_mux_b6/B0_19 ;
  wire  \inst_doa_mux_b6/B0_2 ;
  wire  \inst_doa_mux_b6/B0_20 ;
  wire  \inst_doa_mux_b6/B0_21 ;
  wire  \inst_doa_mux_b6/B0_22 ;
  wire  \inst_doa_mux_b6/B0_23 ;
  wire  \inst_doa_mux_b6/B0_24 ;
  wire  \inst_doa_mux_b6/B0_25 ;
  wire  \inst_doa_mux_b6/B0_26 ;
  wire  \inst_doa_mux_b6/B0_27 ;
  wire  \inst_doa_mux_b6/B0_28 ;
  wire  \inst_doa_mux_b6/B0_29 ;
  wire  \inst_doa_mux_b6/B0_3 ;
  wire  \inst_doa_mux_b6/B0_30 ;
  wire  \inst_doa_mux_b6/B0_31 ;
  wire  \inst_doa_mux_b6/B0_4 ;
  wire  \inst_doa_mux_b6/B0_5 ;
  wire  \inst_doa_mux_b6/B0_6 ;
  wire  \inst_doa_mux_b6/B0_7 ;
  wire  \inst_doa_mux_b6/B0_8 ;
  wire  \inst_doa_mux_b6/B0_9 ;
  wire  \inst_doa_mux_b6/B1_0 ;
  wire  \inst_doa_mux_b6/B1_1 ;
  wire  \inst_doa_mux_b6/B1_10 ;
  wire  \inst_doa_mux_b6/B1_11 ;
  wire  \inst_doa_mux_b6/B1_12 ;
  wire  \inst_doa_mux_b6/B1_13 ;
  wire  \inst_doa_mux_b6/B1_14 ;
  wire  \inst_doa_mux_b6/B1_15 ;
  wire  \inst_doa_mux_b6/B1_2 ;
  wire  \inst_doa_mux_b6/B1_3 ;
  wire  \inst_doa_mux_b6/B1_4 ;
  wire  \inst_doa_mux_b6/B1_5 ;
  wire  \inst_doa_mux_b6/B1_6 ;
  wire  \inst_doa_mux_b6/B1_7 ;
  wire  \inst_doa_mux_b6/B1_8 ;
  wire  \inst_doa_mux_b6/B1_9 ;
  wire  \inst_doa_mux_b6/B2_0 ;
  wire  \inst_doa_mux_b6/B2_1 ;
  wire  \inst_doa_mux_b6/B2_2 ;
  wire  \inst_doa_mux_b6/B2_3 ;
  wire  \inst_doa_mux_b6/B2_4 ;
  wire  \inst_doa_mux_b6/B2_5 ;
  wire  \inst_doa_mux_b6/B2_6 ;
  wire  \inst_doa_mux_b6/B2_7 ;
  wire  \inst_doa_mux_b6/B3_0 ;
  wire  \inst_doa_mux_b6/B3_1 ;
  wire  \inst_doa_mux_b6/B3_2 ;
  wire  \inst_doa_mux_b6/B3_3 ;
  wire  \inst_doa_mux_b6/B4_0 ;
  wire  \inst_doa_mux_b6/B4_1 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire  \inst_doa_mux_b7/B0_10 ;
  wire  \inst_doa_mux_b7/B0_11 ;
  wire  \inst_doa_mux_b7/B0_12 ;
  wire  \inst_doa_mux_b7/B0_13 ;
  wire  \inst_doa_mux_b7/B0_14 ;
  wire  \inst_doa_mux_b7/B0_15 ;
  wire  \inst_doa_mux_b7/B0_16 ;
  wire  \inst_doa_mux_b7/B0_17 ;
  wire  \inst_doa_mux_b7/B0_18 ;
  wire  \inst_doa_mux_b7/B0_19 ;
  wire  \inst_doa_mux_b7/B0_2 ;
  wire  \inst_doa_mux_b7/B0_20 ;
  wire  \inst_doa_mux_b7/B0_21 ;
  wire  \inst_doa_mux_b7/B0_22 ;
  wire  \inst_doa_mux_b7/B0_23 ;
  wire  \inst_doa_mux_b7/B0_24 ;
  wire  \inst_doa_mux_b7/B0_25 ;
  wire  \inst_doa_mux_b7/B0_26 ;
  wire  \inst_doa_mux_b7/B0_27 ;
  wire  \inst_doa_mux_b7/B0_28 ;
  wire  \inst_doa_mux_b7/B0_29 ;
  wire  \inst_doa_mux_b7/B0_3 ;
  wire  \inst_doa_mux_b7/B0_30 ;
  wire  \inst_doa_mux_b7/B0_31 ;
  wire  \inst_doa_mux_b7/B0_4 ;
  wire  \inst_doa_mux_b7/B0_5 ;
  wire  \inst_doa_mux_b7/B0_6 ;
  wire  \inst_doa_mux_b7/B0_7 ;
  wire  \inst_doa_mux_b7/B0_8 ;
  wire  \inst_doa_mux_b7/B0_9 ;
  wire  \inst_doa_mux_b7/B1_0 ;
  wire  \inst_doa_mux_b7/B1_1 ;
  wire  \inst_doa_mux_b7/B1_10 ;
  wire  \inst_doa_mux_b7/B1_11 ;
  wire  \inst_doa_mux_b7/B1_12 ;
  wire  \inst_doa_mux_b7/B1_13 ;
  wire  \inst_doa_mux_b7/B1_14 ;
  wire  \inst_doa_mux_b7/B1_15 ;
  wire  \inst_doa_mux_b7/B1_2 ;
  wire  \inst_doa_mux_b7/B1_3 ;
  wire  \inst_doa_mux_b7/B1_4 ;
  wire  \inst_doa_mux_b7/B1_5 ;
  wire  \inst_doa_mux_b7/B1_6 ;
  wire  \inst_doa_mux_b7/B1_7 ;
  wire  \inst_doa_mux_b7/B1_8 ;
  wire  \inst_doa_mux_b7/B1_9 ;
  wire  \inst_doa_mux_b7/B2_0 ;
  wire  \inst_doa_mux_b7/B2_1 ;
  wire  \inst_doa_mux_b7/B2_2 ;
  wire  \inst_doa_mux_b7/B2_3 ;
  wire  \inst_doa_mux_b7/B2_4 ;
  wire  \inst_doa_mux_b7/B2_5 ;
  wire  \inst_doa_mux_b7/B2_6 ;
  wire  \inst_doa_mux_b7/B2_7 ;
  wire  \inst_doa_mux_b7/B3_0 ;
  wire  \inst_doa_mux_b7/B3_1 ;
  wire  \inst_doa_mux_b7/B3_2 ;
  wire  \inst_doa_mux_b7/B3_3 ;
  wire  \inst_doa_mux_b7/B4_0 ;
  wire  \inst_doa_mux_b7/B4_1 ;
  wire  \inst_doa_mux_b8/B0_0 ;
  wire  \inst_doa_mux_b8/B0_1 ;
  wire  \inst_doa_mux_b8/B0_10 ;
  wire  \inst_doa_mux_b8/B0_11 ;
  wire  \inst_doa_mux_b8/B0_12 ;
  wire  \inst_doa_mux_b8/B0_13 ;
  wire  \inst_doa_mux_b8/B0_14 ;
  wire  \inst_doa_mux_b8/B0_15 ;
  wire  \inst_doa_mux_b8/B0_16 ;
  wire  \inst_doa_mux_b8/B0_17 ;
  wire  \inst_doa_mux_b8/B0_18 ;
  wire  \inst_doa_mux_b8/B0_19 ;
  wire  \inst_doa_mux_b8/B0_2 ;
  wire  \inst_doa_mux_b8/B0_20 ;
  wire  \inst_doa_mux_b8/B0_21 ;
  wire  \inst_doa_mux_b8/B0_22 ;
  wire  \inst_doa_mux_b8/B0_23 ;
  wire  \inst_doa_mux_b8/B0_24 ;
  wire  \inst_doa_mux_b8/B0_25 ;
  wire  \inst_doa_mux_b8/B0_26 ;
  wire  \inst_doa_mux_b8/B0_27 ;
  wire  \inst_doa_mux_b8/B0_28 ;
  wire  \inst_doa_mux_b8/B0_29 ;
  wire  \inst_doa_mux_b8/B0_3 ;
  wire  \inst_doa_mux_b8/B0_30 ;
  wire  \inst_doa_mux_b8/B0_31 ;
  wire  \inst_doa_mux_b8/B0_4 ;
  wire  \inst_doa_mux_b8/B0_5 ;
  wire  \inst_doa_mux_b8/B0_6 ;
  wire  \inst_doa_mux_b8/B0_7 ;
  wire  \inst_doa_mux_b8/B0_8 ;
  wire  \inst_doa_mux_b8/B0_9 ;
  wire  \inst_doa_mux_b8/B1_0 ;
  wire  \inst_doa_mux_b8/B1_1 ;
  wire  \inst_doa_mux_b8/B1_10 ;
  wire  \inst_doa_mux_b8/B1_11 ;
  wire  \inst_doa_mux_b8/B1_12 ;
  wire  \inst_doa_mux_b8/B1_13 ;
  wire  \inst_doa_mux_b8/B1_14 ;
  wire  \inst_doa_mux_b8/B1_15 ;
  wire  \inst_doa_mux_b8/B1_2 ;
  wire  \inst_doa_mux_b8/B1_3 ;
  wire  \inst_doa_mux_b8/B1_4 ;
  wire  \inst_doa_mux_b8/B1_5 ;
  wire  \inst_doa_mux_b8/B1_6 ;
  wire  \inst_doa_mux_b8/B1_7 ;
  wire  \inst_doa_mux_b8/B1_8 ;
  wire  \inst_doa_mux_b8/B1_9 ;
  wire  \inst_doa_mux_b8/B2_0 ;
  wire  \inst_doa_mux_b8/B2_1 ;
  wire  \inst_doa_mux_b8/B2_2 ;
  wire  \inst_doa_mux_b8/B2_3 ;
  wire  \inst_doa_mux_b8/B2_4 ;
  wire  \inst_doa_mux_b8/B2_5 ;
  wire  \inst_doa_mux_b8/B2_6 ;
  wire  \inst_doa_mux_b8/B2_7 ;
  wire  \inst_doa_mux_b8/B3_0 ;
  wire  \inst_doa_mux_b8/B3_1 ;
  wire  \inst_doa_mux_b8/B3_2 ;
  wire  \inst_doa_mux_b8/B3_3 ;
  wire  \inst_doa_mux_b8/B4_0 ;
  wire  \inst_doa_mux_b8/B4_1 ;
  wire \and_Naddra[12]_Naddr_o ;
  wire \and_Naddra[12]_Naddr_o_al_n28 ;
  wire \and_Naddra[12]_Naddr_o_al_n60 ;
  wire \and_Naddra[12]_Naddr_o_al_n92 ;
  wire \and_Naddra[12]_addra_o ;
  wire \and_Naddra[12]_addra_o_al_n108 ;
  wire \and_Naddra[12]_addra_o_al_n44 ;
  wire \and_Naddra[12]_addra_o_al_n76 ;
  wire \and_addra[12]_Naddra_o ;
  wire \and_addra[12]_Naddra_o_al_n100 ;
  wire \and_addra[12]_Naddra_o_al_n36 ;
  wire \and_addra[12]_Naddra_o_al_n68 ;
  wire \and_addra[12]_addra[_o ;
  wire \and_addra[12]_addra[_o_al_n116 ;
  wire \and_addra[12]_addra[_o_al_n52 ;
  wire \and_addra[12]_addra[_o_al_n84 ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i0_008;
  wire inst_doa_i10_000;
  wire inst_doa_i10_001;
  wire inst_doa_i10_002;
  wire inst_doa_i10_003;
  wire inst_doa_i10_004;
  wire inst_doa_i10_005;
  wire inst_doa_i10_006;
  wire inst_doa_i10_007;
  wire inst_doa_i10_008;
  wire inst_doa_i11_000;
  wire inst_doa_i11_001;
  wire inst_doa_i11_002;
  wire inst_doa_i11_003;
  wire inst_doa_i11_004;
  wire inst_doa_i11_005;
  wire inst_doa_i11_006;
  wire inst_doa_i11_007;
  wire inst_doa_i11_008;
  wire inst_doa_i12_000;
  wire inst_doa_i12_001;
  wire inst_doa_i12_002;
  wire inst_doa_i12_003;
  wire inst_doa_i12_004;
  wire inst_doa_i12_005;
  wire inst_doa_i12_006;
  wire inst_doa_i12_007;
  wire inst_doa_i12_008;
  wire inst_doa_i13_000;
  wire inst_doa_i13_001;
  wire inst_doa_i13_002;
  wire inst_doa_i13_003;
  wire inst_doa_i13_004;
  wire inst_doa_i13_005;
  wire inst_doa_i13_006;
  wire inst_doa_i13_007;
  wire inst_doa_i13_008;
  wire inst_doa_i14_000;
  wire inst_doa_i14_001;
  wire inst_doa_i14_002;
  wire inst_doa_i14_003;
  wire inst_doa_i14_004;
  wire inst_doa_i14_005;
  wire inst_doa_i14_006;
  wire inst_doa_i14_007;
  wire inst_doa_i14_008;
  wire inst_doa_i15_000;
  wire inst_doa_i15_001;
  wire inst_doa_i15_002;
  wire inst_doa_i15_003;
  wire inst_doa_i15_004;
  wire inst_doa_i15_005;
  wire inst_doa_i15_006;
  wire inst_doa_i15_007;
  wire inst_doa_i15_008;
  wire inst_doa_i16_000;
  wire inst_doa_i16_001;
  wire inst_doa_i16_002;
  wire inst_doa_i16_003;
  wire inst_doa_i16_004;
  wire inst_doa_i16_005;
  wire inst_doa_i16_006;
  wire inst_doa_i16_007;
  wire inst_doa_i16_008;
  wire inst_doa_i17_000;
  wire inst_doa_i17_001;
  wire inst_doa_i17_002;
  wire inst_doa_i17_003;
  wire inst_doa_i17_004;
  wire inst_doa_i17_005;
  wire inst_doa_i17_006;
  wire inst_doa_i17_007;
  wire inst_doa_i17_008;
  wire inst_doa_i18_000;
  wire inst_doa_i18_001;
  wire inst_doa_i18_002;
  wire inst_doa_i18_003;
  wire inst_doa_i18_004;
  wire inst_doa_i18_005;
  wire inst_doa_i18_006;
  wire inst_doa_i18_007;
  wire inst_doa_i18_008;
  wire inst_doa_i19_000;
  wire inst_doa_i19_001;
  wire inst_doa_i19_002;
  wire inst_doa_i19_003;
  wire inst_doa_i19_004;
  wire inst_doa_i19_005;
  wire inst_doa_i19_006;
  wire inst_doa_i19_007;
  wire inst_doa_i19_008;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i1_008;
  wire inst_doa_i20_000;
  wire inst_doa_i20_001;
  wire inst_doa_i20_002;
  wire inst_doa_i20_003;
  wire inst_doa_i20_004;
  wire inst_doa_i20_005;
  wire inst_doa_i20_006;
  wire inst_doa_i20_007;
  wire inst_doa_i20_008;
  wire inst_doa_i21_000;
  wire inst_doa_i21_001;
  wire inst_doa_i21_002;
  wire inst_doa_i21_003;
  wire inst_doa_i21_004;
  wire inst_doa_i21_005;
  wire inst_doa_i21_006;
  wire inst_doa_i21_007;
  wire inst_doa_i21_008;
  wire inst_doa_i22_000;
  wire inst_doa_i22_001;
  wire inst_doa_i22_002;
  wire inst_doa_i22_003;
  wire inst_doa_i22_004;
  wire inst_doa_i22_005;
  wire inst_doa_i22_006;
  wire inst_doa_i22_007;
  wire inst_doa_i22_008;
  wire inst_doa_i23_000;
  wire inst_doa_i23_001;
  wire inst_doa_i23_002;
  wire inst_doa_i23_003;
  wire inst_doa_i23_004;
  wire inst_doa_i23_005;
  wire inst_doa_i23_006;
  wire inst_doa_i23_007;
  wire inst_doa_i23_008;
  wire inst_doa_i24_000;
  wire inst_doa_i24_001;
  wire inst_doa_i24_002;
  wire inst_doa_i24_003;
  wire inst_doa_i24_004;
  wire inst_doa_i24_005;
  wire inst_doa_i24_006;
  wire inst_doa_i24_007;
  wire inst_doa_i24_008;
  wire inst_doa_i25_000;
  wire inst_doa_i25_001;
  wire inst_doa_i25_002;
  wire inst_doa_i25_003;
  wire inst_doa_i25_004;
  wire inst_doa_i25_005;
  wire inst_doa_i25_006;
  wire inst_doa_i25_007;
  wire inst_doa_i25_008;
  wire inst_doa_i26_000;
  wire inst_doa_i26_001;
  wire inst_doa_i26_002;
  wire inst_doa_i26_003;
  wire inst_doa_i26_004;
  wire inst_doa_i26_005;
  wire inst_doa_i26_006;
  wire inst_doa_i26_007;
  wire inst_doa_i26_008;
  wire inst_doa_i27_000;
  wire inst_doa_i27_001;
  wire inst_doa_i27_002;
  wire inst_doa_i27_003;
  wire inst_doa_i27_004;
  wire inst_doa_i27_005;
  wire inst_doa_i27_006;
  wire inst_doa_i27_007;
  wire inst_doa_i27_008;
  wire inst_doa_i28_000;
  wire inst_doa_i28_001;
  wire inst_doa_i28_002;
  wire inst_doa_i28_003;
  wire inst_doa_i28_004;
  wire inst_doa_i28_005;
  wire inst_doa_i28_006;
  wire inst_doa_i28_007;
  wire inst_doa_i28_008;
  wire inst_doa_i29_000;
  wire inst_doa_i29_001;
  wire inst_doa_i29_002;
  wire inst_doa_i29_003;
  wire inst_doa_i29_004;
  wire inst_doa_i29_005;
  wire inst_doa_i29_006;
  wire inst_doa_i29_007;
  wire inst_doa_i29_008;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;
  wire inst_doa_i2_008;
  wire inst_doa_i30_000;
  wire inst_doa_i30_001;
  wire inst_doa_i30_002;
  wire inst_doa_i30_003;
  wire inst_doa_i30_004;
  wire inst_doa_i30_005;
  wire inst_doa_i30_006;
  wire inst_doa_i30_007;
  wire inst_doa_i30_008;
  wire inst_doa_i31_000;
  wire inst_doa_i31_001;
  wire inst_doa_i31_002;
  wire inst_doa_i31_003;
  wire inst_doa_i31_004;
  wire inst_doa_i31_005;
  wire inst_doa_i31_006;
  wire inst_doa_i31_007;
  wire inst_doa_i31_008;
  wire inst_doa_i32_000;
  wire inst_doa_i32_001;
  wire inst_doa_i32_002;
  wire inst_doa_i32_003;
  wire inst_doa_i32_004;
  wire inst_doa_i32_005;
  wire inst_doa_i32_006;
  wire inst_doa_i32_007;
  wire inst_doa_i32_008;
  wire inst_doa_i33_000;
  wire inst_doa_i33_001;
  wire inst_doa_i33_002;
  wire inst_doa_i33_003;
  wire inst_doa_i33_004;
  wire inst_doa_i33_005;
  wire inst_doa_i33_006;
  wire inst_doa_i33_007;
  wire inst_doa_i33_008;
  wire inst_doa_i34_000;
  wire inst_doa_i34_001;
  wire inst_doa_i34_002;
  wire inst_doa_i34_003;
  wire inst_doa_i34_004;
  wire inst_doa_i34_005;
  wire inst_doa_i34_006;
  wire inst_doa_i34_007;
  wire inst_doa_i34_008;
  wire inst_doa_i35_000;
  wire inst_doa_i35_001;
  wire inst_doa_i35_002;
  wire inst_doa_i35_003;
  wire inst_doa_i35_004;
  wire inst_doa_i35_005;
  wire inst_doa_i35_006;
  wire inst_doa_i35_007;
  wire inst_doa_i35_008;
  wire inst_doa_i36_000;
  wire inst_doa_i36_001;
  wire inst_doa_i36_002;
  wire inst_doa_i36_003;
  wire inst_doa_i36_004;
  wire inst_doa_i36_005;
  wire inst_doa_i36_006;
  wire inst_doa_i36_007;
  wire inst_doa_i36_008;
  wire inst_doa_i37_000;
  wire inst_doa_i37_001;
  wire inst_doa_i37_002;
  wire inst_doa_i37_003;
  wire inst_doa_i37_004;
  wire inst_doa_i37_005;
  wire inst_doa_i37_006;
  wire inst_doa_i37_007;
  wire inst_doa_i37_008;
  wire inst_doa_i38_000;
  wire inst_doa_i38_001;
  wire inst_doa_i38_002;
  wire inst_doa_i38_003;
  wire inst_doa_i38_004;
  wire inst_doa_i38_005;
  wire inst_doa_i38_006;
  wire inst_doa_i38_007;
  wire inst_doa_i38_008;
  wire inst_doa_i39_000;
  wire inst_doa_i39_001;
  wire inst_doa_i39_002;
  wire inst_doa_i39_003;
  wire inst_doa_i39_004;
  wire inst_doa_i39_005;
  wire inst_doa_i39_006;
  wire inst_doa_i39_007;
  wire inst_doa_i39_008;
  wire inst_doa_i3_000;
  wire inst_doa_i3_001;
  wire inst_doa_i3_002;
  wire inst_doa_i3_003;
  wire inst_doa_i3_004;
  wire inst_doa_i3_005;
  wire inst_doa_i3_006;
  wire inst_doa_i3_007;
  wire inst_doa_i3_008;
  wire inst_doa_i40_000;
  wire inst_doa_i40_001;
  wire inst_doa_i40_002;
  wire inst_doa_i40_003;
  wire inst_doa_i40_004;
  wire inst_doa_i40_005;
  wire inst_doa_i40_006;
  wire inst_doa_i40_007;
  wire inst_doa_i40_008;
  wire inst_doa_i41_000;
  wire inst_doa_i41_001;
  wire inst_doa_i41_002;
  wire inst_doa_i41_003;
  wire inst_doa_i41_004;
  wire inst_doa_i41_005;
  wire inst_doa_i41_006;
  wire inst_doa_i41_007;
  wire inst_doa_i41_008;
  wire inst_doa_i42_000;
  wire inst_doa_i42_001;
  wire inst_doa_i42_002;
  wire inst_doa_i42_003;
  wire inst_doa_i42_004;
  wire inst_doa_i42_005;
  wire inst_doa_i42_006;
  wire inst_doa_i42_007;
  wire inst_doa_i42_008;
  wire inst_doa_i43_000;
  wire inst_doa_i43_001;
  wire inst_doa_i43_002;
  wire inst_doa_i43_003;
  wire inst_doa_i43_004;
  wire inst_doa_i43_005;
  wire inst_doa_i43_006;
  wire inst_doa_i43_007;
  wire inst_doa_i43_008;
  wire inst_doa_i44_000;
  wire inst_doa_i44_001;
  wire inst_doa_i44_002;
  wire inst_doa_i44_003;
  wire inst_doa_i44_004;
  wire inst_doa_i44_005;
  wire inst_doa_i44_006;
  wire inst_doa_i44_007;
  wire inst_doa_i44_008;
  wire inst_doa_i45_000;
  wire inst_doa_i45_001;
  wire inst_doa_i45_002;
  wire inst_doa_i45_003;
  wire inst_doa_i45_004;
  wire inst_doa_i45_005;
  wire inst_doa_i45_006;
  wire inst_doa_i45_007;
  wire inst_doa_i45_008;
  wire inst_doa_i46_000;
  wire inst_doa_i46_001;
  wire inst_doa_i46_002;
  wire inst_doa_i46_003;
  wire inst_doa_i46_004;
  wire inst_doa_i46_005;
  wire inst_doa_i46_006;
  wire inst_doa_i46_007;
  wire inst_doa_i46_008;
  wire inst_doa_i47_000;
  wire inst_doa_i47_001;
  wire inst_doa_i47_002;
  wire inst_doa_i47_003;
  wire inst_doa_i47_004;
  wire inst_doa_i47_005;
  wire inst_doa_i47_006;
  wire inst_doa_i47_007;
  wire inst_doa_i47_008;
  wire inst_doa_i48_000;
  wire inst_doa_i48_001;
  wire inst_doa_i48_002;
  wire inst_doa_i48_003;
  wire inst_doa_i48_004;
  wire inst_doa_i48_005;
  wire inst_doa_i48_006;
  wire inst_doa_i48_007;
  wire inst_doa_i48_008;
  wire inst_doa_i49_000;
  wire inst_doa_i49_001;
  wire inst_doa_i49_002;
  wire inst_doa_i49_003;
  wire inst_doa_i49_004;
  wire inst_doa_i49_005;
  wire inst_doa_i49_006;
  wire inst_doa_i49_007;
  wire inst_doa_i49_008;
  wire inst_doa_i4_000;
  wire inst_doa_i4_001;
  wire inst_doa_i4_002;
  wire inst_doa_i4_003;
  wire inst_doa_i4_004;
  wire inst_doa_i4_005;
  wire inst_doa_i4_006;
  wire inst_doa_i4_007;
  wire inst_doa_i4_008;
  wire inst_doa_i50_000;
  wire inst_doa_i50_001;
  wire inst_doa_i50_002;
  wire inst_doa_i50_003;
  wire inst_doa_i50_004;
  wire inst_doa_i50_005;
  wire inst_doa_i50_006;
  wire inst_doa_i50_007;
  wire inst_doa_i50_008;
  wire inst_doa_i51_000;
  wire inst_doa_i51_001;
  wire inst_doa_i51_002;
  wire inst_doa_i51_003;
  wire inst_doa_i51_004;
  wire inst_doa_i51_005;
  wire inst_doa_i51_006;
  wire inst_doa_i51_007;
  wire inst_doa_i51_008;
  wire inst_doa_i52_000;
  wire inst_doa_i52_001;
  wire inst_doa_i52_002;
  wire inst_doa_i52_003;
  wire inst_doa_i52_004;
  wire inst_doa_i52_005;
  wire inst_doa_i52_006;
  wire inst_doa_i52_007;
  wire inst_doa_i52_008;
  wire inst_doa_i53_000;
  wire inst_doa_i53_001;
  wire inst_doa_i53_002;
  wire inst_doa_i53_003;
  wire inst_doa_i53_004;
  wire inst_doa_i53_005;
  wire inst_doa_i53_006;
  wire inst_doa_i53_007;
  wire inst_doa_i53_008;
  wire inst_doa_i54_000;
  wire inst_doa_i54_001;
  wire inst_doa_i54_002;
  wire inst_doa_i54_003;
  wire inst_doa_i54_004;
  wire inst_doa_i54_005;
  wire inst_doa_i54_006;
  wire inst_doa_i54_007;
  wire inst_doa_i54_008;
  wire inst_doa_i55_000;
  wire inst_doa_i55_001;
  wire inst_doa_i55_002;
  wire inst_doa_i55_003;
  wire inst_doa_i55_004;
  wire inst_doa_i55_005;
  wire inst_doa_i55_006;
  wire inst_doa_i55_007;
  wire inst_doa_i55_008;
  wire inst_doa_i56_000;
  wire inst_doa_i56_001;
  wire inst_doa_i56_002;
  wire inst_doa_i56_003;
  wire inst_doa_i56_004;
  wire inst_doa_i56_005;
  wire inst_doa_i56_006;
  wire inst_doa_i56_007;
  wire inst_doa_i56_008;
  wire inst_doa_i57_000;
  wire inst_doa_i57_001;
  wire inst_doa_i57_002;
  wire inst_doa_i57_003;
  wire inst_doa_i57_004;
  wire inst_doa_i57_005;
  wire inst_doa_i57_006;
  wire inst_doa_i57_007;
  wire inst_doa_i57_008;
  wire inst_doa_i58_000;
  wire inst_doa_i58_001;
  wire inst_doa_i58_002;
  wire inst_doa_i58_003;
  wire inst_doa_i58_004;
  wire inst_doa_i58_005;
  wire inst_doa_i58_006;
  wire inst_doa_i58_007;
  wire inst_doa_i58_008;
  wire inst_doa_i59_000;
  wire inst_doa_i59_001;
  wire inst_doa_i59_002;
  wire inst_doa_i59_003;
  wire inst_doa_i59_004;
  wire inst_doa_i59_005;
  wire inst_doa_i59_006;
  wire inst_doa_i59_007;
  wire inst_doa_i59_008;
  wire inst_doa_i5_000;
  wire inst_doa_i5_001;
  wire inst_doa_i5_002;
  wire inst_doa_i5_003;
  wire inst_doa_i5_004;
  wire inst_doa_i5_005;
  wire inst_doa_i5_006;
  wire inst_doa_i5_007;
  wire inst_doa_i5_008;
  wire inst_doa_i60_000;
  wire inst_doa_i60_001;
  wire inst_doa_i60_002;
  wire inst_doa_i60_003;
  wire inst_doa_i60_004;
  wire inst_doa_i60_005;
  wire inst_doa_i60_006;
  wire inst_doa_i60_007;
  wire inst_doa_i60_008;
  wire inst_doa_i61_000;
  wire inst_doa_i61_001;
  wire inst_doa_i61_002;
  wire inst_doa_i61_003;
  wire inst_doa_i61_004;
  wire inst_doa_i61_005;
  wire inst_doa_i61_006;
  wire inst_doa_i61_007;
  wire inst_doa_i61_008;
  wire inst_doa_i62_000;
  wire inst_doa_i62_001;
  wire inst_doa_i62_002;
  wire inst_doa_i62_003;
  wire inst_doa_i62_004;
  wire inst_doa_i62_005;
  wire inst_doa_i62_006;
  wire inst_doa_i62_007;
  wire inst_doa_i62_008;
  wire inst_doa_i63_000;
  wire inst_doa_i63_001;
  wire inst_doa_i63_002;
  wire inst_doa_i63_003;
  wire inst_doa_i63_004;
  wire inst_doa_i63_005;
  wire inst_doa_i63_006;
  wire inst_doa_i63_007;
  wire inst_doa_i63_008;
  wire inst_doa_i6_000;
  wire inst_doa_i6_001;
  wire inst_doa_i6_002;
  wire inst_doa_i6_003;
  wire inst_doa_i6_004;
  wire inst_doa_i6_005;
  wire inst_doa_i6_006;
  wire inst_doa_i6_007;
  wire inst_doa_i6_008;
  wire inst_doa_i7_000;
  wire inst_doa_i7_001;
  wire inst_doa_i7_002;
  wire inst_doa_i7_003;
  wire inst_doa_i7_004;
  wire inst_doa_i7_005;
  wire inst_doa_i7_006;
  wire inst_doa_i7_007;
  wire inst_doa_i7_008;
  wire inst_doa_i8_000;
  wire inst_doa_i8_001;
  wire inst_doa_i8_002;
  wire inst_doa_i8_003;
  wire inst_doa_i8_004;
  wire inst_doa_i8_005;
  wire inst_doa_i8_006;
  wire inst_doa_i8_007;
  wire inst_doa_i8_008;
  wire inst_doa_i9_000;
  wire inst_doa_i9_001;
  wire inst_doa_i9_002;
  wire inst_doa_i9_003;
  wire inst_doa_i9_004;
  wire inst_doa_i9_005;
  wire inst_doa_i9_006;
  wire inst_doa_i9_007;
  wire inst_doa_i9_008;

  reg_sr_as_w1 addra_pipe_b0 (
    .clk(clka),
    .d(addra[10]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[0]));
  reg_sr_as_w1 addra_pipe_b1 (
    .clk(clka),
    .d(addra[11]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[1]));
  reg_sr_as_w1 addra_pipe_b2 (
    .clk(clka),
    .d(addra[12]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[2]));
  reg_sr_as_w1 addra_pipe_b3 (
    .clk(clka),
    .d(addra[13]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[3]));
  reg_sr_as_w1 addra_pipe_b4 (
    .clk(clka),
    .d(addra[14]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[4]));
  reg_sr_as_w1 addra_pipe_b5 (
    .clk(clka),
    .d(addra[15]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[5]));
  and \and_Naddra[12]_Naddr  (\and_Naddra[12]_Naddr_o , ~addra[12], ~addra[13], ~addra[14], ~addra[15]);
  and \and_Naddra[12]_Naddr_al_u28  (\and_Naddra[12]_Naddr_o_al_n28 , ~addra[12], ~addra[13], addra[14], ~addra[15]);
  and \and_Naddra[12]_Naddr_al_u60  (\and_Naddra[12]_Naddr_o_al_n60 , ~addra[12], ~addra[13], ~addra[14], addra[15]);
  and \and_Naddra[12]_Naddr_al_u92  (\and_Naddra[12]_Naddr_o_al_n92 , ~addra[12], ~addra[13], addra[14], addra[15]);
  and \and_Naddra[12]_addra  (\and_Naddra[12]_addra_o , ~addra[12], addra[13], ~addra[14], ~addra[15]);
  and \and_Naddra[12]_addra_al_u108  (\and_Naddra[12]_addra_o_al_n108 , ~addra[12], addra[13], addra[14], addra[15]);
  and \and_Naddra[12]_addra_al_u44  (\and_Naddra[12]_addra_o_al_n44 , ~addra[12], addra[13], addra[14], ~addra[15]);
  and \and_Naddra[12]_addra_al_u76  (\and_Naddra[12]_addra_o_al_n76 , ~addra[12], addra[13], ~addra[14], addra[15]);
  and \and_addra[12]_Naddra  (\and_addra[12]_Naddra_o , addra[12], ~addra[13], ~addra[14], ~addra[15]);
  and \and_addra[12]_Naddra_al_u100  (\and_addra[12]_Naddra_o_al_n100 , addra[12], ~addra[13], addra[14], addra[15]);
  and \and_addra[12]_Naddra_al_u36  (\and_addra[12]_Naddra_o_al_n36 , addra[12], ~addra[13], addra[14], ~addra[15]);
  and \and_addra[12]_Naddra_al_u68  (\and_addra[12]_Naddra_o_al_n68 , addra[12], ~addra[13], ~addra[14], addra[15]);
  and \and_addra[12]_addra[  (\and_addra[12]_addra[_o , addra[12], addra[13], ~addra[14], ~addra[15]);
  and \and_addra[12]_addra[_al_u116  (\and_addra[12]_addra[_o_al_n116 , addra[12], addra[13], addra[14], addra[15]);
  and \and_addra[12]_addra[_al_u52  (\and_addra[12]_addra[_o_al_n52 , addra[12], addra[13], addra[14], ~addra[15]);
  and \and_addra[12]_addra[_al_u84  (\and_addra[12]_addra[_o_al_n84 , addra[12], addra[13], ~addra[14], addra[15]);
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hF6FFFFF7F6F6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFF6F7F7FFFFF6F6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7B6FFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFF66D2424246C6DB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_000000_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_008,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFF6D1B6DB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFB6B6FFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFF2464FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFAE6D6D6DB6FFFFFFFFFFFFFFFFFFB66DB6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFF6B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hB6FFFFFFB6FFFFFFF7FFFFFFFFFFFFFFFFFFF6F7FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFF246DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFAE25656E651C65AEF7FFFFFFFFFFF7DBD31C25AEF7FFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFB6F6FFFFFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFAEB6F7B6F7FFFFF7B6F6FFF7F6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFF6D6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFB624656666666E652525656DB6FFF71C9393D31C1C65B6FFFFFFFFFFFFFF),
    .INIT_1E(256'hF6ADFFFFFFF7FFF6F6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hF6FFF7F7FFFFF7FFF7F6B6F6FFFFFFFFFFFFFFFFF6FFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_001024_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_008,inst_doa_i1_007,inst_doa_i1_006,inst_doa_i1_005,inst_doa_i1_004,inst_doa_i1_003,inst_doa_i1_002,inst_doa_i1_001,inst_doa_i1_000}));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFCF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFE79FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFC7FBCFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFF03FDE7FFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFF24FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFF25656566666666656565251C8AD36565251C8B931C1C24AEFFFFFFFFFFFF),
    .INIT_06(256'hFFF6FFFFF6AEF6F7F7FFADFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hB6B6FFFFB6F6FFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6FFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFF6DFFFFB6ADADB6B6F6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFF6D1C656566656566656565656565D3D36566651DD38B1D1D1C6DFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFB6FFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFF7FFB6B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFB6AD6464DAD21B2364646DADB6B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hF71C2565651C8A42D4656666656565661C8B65AE651DD48B1D1C246DFFFFFFFF),
    .INIT_16(256'hFFFFFFB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6F6FFFFFF),
    .INIT_17(256'hFFF6FFFFFFFFB6B6FFFFFFFFFFB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h6C241BDB89481B6464646464646CADB6B6B6F6FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6),
    .INIT_1D(256'h651C6565D48A8A8A418A1C66AE661D1D1D1CD365AE651DD48B251C25AEFFFFFF),
    .INIT_1E(256'hFFB66DB6F6FFB6B6ADB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6F7F6F6FFFF),
    .INIT_1F(256'hF66DFFFFFFFFFF6DFFB6B6B66DADF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_002048_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i2_008,inst_doa_i2_007,inst_doa_i2_006,inst_doa_i2_005,inst_doa_i2_004,inst_doa_i2_003,inst_doa_i2_002,inst_doa_i2_001,inst_doa_i2_000}));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFF600FEF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFC007F79FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFE807FCBDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFD81FFF5EFFFFFFFFFFFFFFFFFFFFFFFFFFE03BFFFFFFFFFFF),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFB6B6B6AD6D6D6D6D6D6D6DB6B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'h64646464641B6364646464646464646C6DAD6DADB6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF66C24),
    .INIT_05(256'hD3651C938A8A8A8A8B8A41D3656E66651D1D1CD365AE651DD4D31D1C65246DB6),
    .INIT_06(256'hF6FFB6FFFFB6B6B6F6B6B6B6B6B6FFFFFFFFFFFFFFFFFFFFFFF6B6FFFFFFFFF7),
    .INIT_07(256'hB6ADFFFFFFFFFFB6FFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hB66D6D6D6D6D6D6D6D6D6D6D6D6424246DADB6FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h646464646464646464646464646464646464646C646DB6FFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h25AEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAD242364),
    .INIT_0D(256'h1C1DD38A8A8A8A8A8A8B8B8A8A256665651D1D1CD365AE6525D4D41D1C651C65),
    .INIT_0E(256'hFFFFFFFFFFFFFFF6FFFFF6F6FFFFFFB6F6FFFFFFFFFFFFFFFFFFFFFFFFFFFF65),
    .INIT_0F(256'hB6B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFFFFFFFFFFFFB6B6AE),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hB5B5B6B6B6B6ADAD6D6D6D6D6D6C2424246C6D6DB6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6B6),
    .INIT_13(256'h64646464646464646464646464646464646464646C64646DFFFFFFFFFFFFFFFF),
    .INIT_14(256'h6D2465B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6D23236464),
    .INIT_15(256'h1DD48B8A8A8A8AD3D41C1D65651C65651D25DCDC1CD36EAE6525D31C1D1D6565),
    .INIT_16(256'hF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFB665D3),
    .INIT_17(256'hFFB6FFFFAEB6FFFFFFFFFFFFB6FFFFFFFFFFF6F6B6F6FFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hB6F6B6B66D2424DBDBDBDBDBDBDB1B1B1BDB246DB6B6B6FFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6B6B6),
    .INIT_1B(256'h6D6D6464646464646464646464646464646464646464646464B6FFFFFFFFFFFF),
    .INIT_1C(256'h656E6524AEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF64241B646464),
    .INIT_1D(256'h1C8B8A8A8B8AD31C65656566666E65656565251CDC1CD366AE6525D31D1D1D65),
    .INIT_1E(256'hF7B6FFFFFFFFFFFFFFB6B6FFFFFFFFFFFFFFFFFFB6F7FFFFFFFFFFB6651CDC1C),
    .INIT_1F(256'hFFF6FFFFFFFFFFFFFFF6FFB6ADFFFFFFFFFFF6F6FFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_003072_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i3_008,inst_doa_i3_007,inst_doa_i3_006,inst_doa_i3_005,inst_doa_i3_004,inst_doa_i3_003,inst_doa_i3_002,inst_doa_i3_001,inst_doa_i3_000}));
  // address_offset=4096;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFBD03FFFCF7FFFFFFFFFFFFFFFFFFFFFFFFE0037FFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFEC07FFFF7BFFFFFFFFFFFFFFFFFFFFFFFF8001FFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFBFF003FFFF9FFFFFFF7FFFFFFFFFFFFFFFFE00032FFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFF61F81FFFFFEFFF7FFE7FFFFFFFFFFFFFFFF8000EFF7FFFFFFFFF),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFB665DB924949929292DBDBDBDB241CDB2424246DB6F6B6B6FFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6FEF6B6FE),
    .INIT_03(256'hAD6C6C6464646C6C6C6464646464646464646464646464646424ADFFFFFFFFFF),
    .INIT_04(256'h65666E652565FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2423231B6C64AD),
    .INIT_05(256'hD38A8A8B8BD32566666665656565656565656E66651CD4D36EAE661DD31D1D65),
    .INIT_06(256'hFFF6FFFFFFFFFFFFF6ADB6B6FFFFFFFFFFFFB6AE6DB6F7F765DC1C1D6565D41C),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFB6B6FFFFFFFFFFFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h249249494992929292929292DBDB921C6C24242424246DB6B6ADFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6FEB6B6F6B6),
    .INIT_0B(256'hADACAC6C64646CADADADAC6464646464646464646464646464646464FFFFFFFF),
    .INIT_0C(256'h65656E66662524FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF641B641B6463ADB5),
    .INIT_0D(256'h8B8A8BD3D31C656565666EAEAEAEAE6E656565656E6E661CDC6566661CD41D1D),
    .INIT_0E(256'hFFFFFFFFB6FFFFFFFFB6FFFFFFFFFFFFF72424656D656D65651C1CDC251DD3D4),
    .INIT_0F(256'hF6FFFFFFFFFFFFFFFFFFB6FFFFFFB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h00499292929292919292D2DA92DB2464DBDB1BDB24242424B6F66DB6FFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6B6B6B6B62449),
    .INIT_13(256'hADAD6C6463ADADADAC6464646464646464646464646464646464646464B6FFFF),
    .INIT_14(256'h1D6566AE6665651CF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFB592641B64646CF5AD),
    .INIT_15(256'h8B8A8B8BD3D41C1D656565666EAEB7B7B7AEAEAE6E6E6EAE65DCD425661C1C1D),
    .INIT_16(256'hFFF7FFFFFFB6FFFFFFFFFFFFFFFFFFFFAEDC6565656565656566651CD3D3D3D3),
    .INIT_17(256'hF6FFFFF6FFFFFFFFFFF7AEFFF7FFB6B6FFFFFFFFF6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h49924949494992DADBDB92DA646D64DB246D6D241B242424DB24B66DB6FFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB5B6B6ADB56D920049),
    .INIT_1B(256'hAD6C1B236C6C641B1A1B6464646464646464646464646464646464646464F6FF),
    .INIT_1C(256'h1D25656EAE6E6E6DDCF7FFFFFFFFFFFFFFFFFFFFFFFFFFDBDB231B641BF6ADAC),
    .INIT_1D(256'h8A8AD41C1C1C1C1D6565656565656565AEAEB7B7AEAEAEAEAEAE25D31C651C1D),
    .INIT_1E(256'hF6B6F6FFFFB66DFFFFF6F6F6FFFFFFF7D36565D38A8BD41D656525651C8AD38B),
    .INIT_1F(256'hFFF7F6FFF6FFFFFFFFB6AEFFFFB6B6F6B6B6FFF6ADF6FFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_004096_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i4_008,inst_doa_i4_007,inst_doa_i4_006,inst_doa_i4_005,inst_doa_i4_004,inst_doa_i4_003,inst_doa_i4_002,inst_doa_i4_001,inst_doa_i4_000}));
  // address_offset=5120;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFF60783FFFFFF3FFFFFEFFF9FFFFFFFFFFFFF0003FFF9FFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFEC000FFFFFFFCEFFFFCFFA3FFFFFFFFFFFFC010F7FF9FFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFE80007FFFFFFE67FFFDFF0FFFFFFFFFFFFF8061FFFFF7FFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFD800F7FFFFFFF73FFFD7F1DFFFFFFFFFFFF0187FFFDFBFFFFFFFF),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h49494992DADBDBDBD29224AD6D241B646D6D6C64242424646DDBDBB56D6DFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAD6D6D6D6D2300004949),
    .INIT_03(256'h6C1B1B231BD2D21B646C646464646464646464646464646464646464646464F6),
    .INIT_04(256'h1D1C1D656EAE6E6EAE1CF7FFFFFFFFFFFFFFFFFFFFFF6D91241B1B1BACB56CAC),
    .INIT_05(256'h8BD41D65666665656565656565656565656565AEAEAEAEAEAEAEAF66D3D41D1C),
    .INIT_06(256'hF7FFFFFFB6B6B6FFFFFFFFFFFFFFFF25D4661C428B8A42418B1C1C1C1C8B8B8B),
    .INIT_07(256'hFFFFFFF7F6FFFFFFB6B6F7FFFFFFB6B6FFFFFFFFFFF6FFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h4992DB23DBDBD2921B6DB66CDB246D6D6D6D646D6D6D6DB524DBDB246D6D6DFF),
    .INIT_0A(256'hF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6646D6D6DDB0049494949),
    .INIT_0B(256'h1BD21BD248DA6CAD64236464646C646464646464646464646464646464646464),
    .INIT_0C(256'h1D1D1CDC6566AE6E6EAE1CF7FFFFFFFFFFFFFFFFFFFFDBD21B1A631BADAC646C),
    .INIT_0D(256'h1C65656565666EAE656565666EAE6565656EAEAE6565AEAE6EAEAEF7B71C8BDC),
    .INIT_0E(256'hF6F7FFFFF7FFFFFFFFFFFFFFFFFFB78A1D65D38A8B8B8B8B8A8BD3D3D38B8BD3),
    .INIT_0F(256'hFFFFFFF6F6FFFFFFB6B6FFFFFFFFF6F6FFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hDB241BDBDA92DB6DB66D231B6C6D6C6D6D6D6D6D6C6DB51B246D6D24DB6D6D6D),
    .INIT_12(256'h6CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE2424646D92004949000092),
    .INIT_13(256'hDAD292401BADAD1B1B64ADADAC64646464646464646464646464646464646464),
    .INIT_14(256'hDC1D1DD3D46566AF6EAEAE1CF7FFFFFFFFFFFFFFFFB6921B1B1B1B63AD646464),
    .INIT_15(256'hD4656665666565AEAE6E656565AEAEAE6E6565AEB7AE656DAE6E6565AFF7658A),
    .INIT_16(256'hF6F6FFFFFFFFFFFFFFFFFFFFFFFF258B65D4418A8B8A8BD3D38B8B8BD4D4D3D3),
    .INIT_17(256'hFFF7F6F6FFF6FFFFFFFFF6B6FFFFFFF6FFFFF6F6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h24DBDBDAD224B5B5241B646D6D6DAD6DADB66D646D6DDB24AD6D6D6464DA246D),
    .INIT_1A(256'h246DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF24242424920049000091DB24),
    .INIT_1B(256'h92910023AD64D21A6CAD6C646464AD6C64646464646464646464646464646464),
    .INIT_1C(256'hD31C251C93DC6566AF6EAEB61CF7FFFFFFFFFFFFFF6C911BDA1B1A6464236C1B),
    .INIT_1D(256'hD41C666665666565AEF7AE6E65656EAEB7AEAE656DAEB66D6565AE651D6EB766),
    .INIT_1E(256'hF6F6FFFFFFFFFFFFB6FFFFFFFFB7411C1C8BD3D4D4D4D38B8BD38B8A1C651D65),
    .INIT_1F(256'hFFFFF6F6F6FFFFFFFFFFF6B6F6FFF6F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_005120_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i5_008,inst_doa_i5_007,inst_doa_i5_006,inst_doa_i5_005,inst_doa_i5_004,inst_doa_i5_003,inst_doa_i5_002,inst_doa_i5_001,inst_doa_i5_000}));
  // address_offset=6144;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFDF81FFFFFFFFFB9FFF95E1BFFFFFFFFFFF6060EFFFBF9FFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFBFFFFFFFFFFFEDDFFFBFEB3FFFFFFFFFFEC183DFFF7F8F7FFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFF6E7FFABDA67FFFFFDFFFE87277FFEFFE1BFFFFFF),
    .INITP_03(256'hFFFFFFFFFFDFFFFFFFFFFFFDBF7FF2BF8C37FFFFDFFFD0C9EFFFDFFFFDFFFFFF),
    .INIT_00(256'h2424FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hDBDBD2DB6DB66DDB246D6D6DADB5ADB6B66D246D6DDB24B56D6D6C6D64DB9224),
    .INIT_02(256'h6423B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6DDB2424D200490000DB2424DB),
    .INIT_03(256'hD2D2D2AD24481B6CAD64236464ADAD64646464646C6464646464646464646463),
    .INIT_04(256'h66D31C251DD3D46566AF6DB6AE1CF7FFFFFFFFFFFFDBD21BDA1BDA64636464D2),
    .INIT_05(256'h661C25AEAE65656565AEF7AEAE6565656EB7F7B6AE65AEB6AE65256EAE1C1DAE),
    .INIT_06(256'hFFFFFFFFFFFFFFFFF6FFFFFFFF1C4A1D1C65651D1CD4D38BD3D4D41C1D656565),
    .INIT_07(256'hF6F6F7F6F6F7FFFFB6FFFFF6B6F6F6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h24236DB6DB6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hDB9224B6B524DB246DAD6DB5B6B6B6B66D246D6C9224B6AD6D6D64AD24DBDB92),
    .INIT_0A(256'h232364FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6DB2424DB490000922424DBDBDB),
    .INIT_0B(256'h64D2642340D2646C1B1B6363ADAD64636C64646C64646C6C6464646464646464),
    .INIT_0C(256'h6625D31C6525D31C6566AE6EB6AE1CF7FFFFFFFFB6891B1B1A1B1B641B6423D2),
    .INIT_0D(256'h6E6E1C65AEAE656E6E65AEB7AEAE65656565AEB7F7AE6E6DAEAE6D1C65AE25DC),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFF6ED32566AEAE65651C1C1C1D1D1C656565656565),
    .INIT_0F(256'hF7F7FFF6F6F7FFB6B6FFFFFFADF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h49DBDB1B24DB6CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hDB6DB66CDB236CADB5ADB6B6B6B6B524246D249224B5B56D6D6D6DAD24232492),
    .INIT_12(256'h641BDBB5FFFFFFFFFFFFFFFFFFFFFFFFFFFF23DB24DB890000242424DBDB24DA),
    .INIT_13(256'h64D21B89892364DAD21B1AADAD1B636C6464642364AC6C6C6C646464646C646C),
    .INIT_14(256'hD4651CD31D651DD3DC6566AEAEB7AE24FFFFFFFF64891BDA1BD21B641B64DA23),
    .INIT_15(256'h65AEAE6565AEB76E6EAE65AEAEAEAEAE65656565AEF7AEAE6D6E6EAE1C1C6E25),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFF7651C65AEB6AE66656565656566651D666666656566),
    .INIT_17(256'hFFF7F7F6FFFFFFFFFFFFFFFFF6F6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h236424246C24DB6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hB56D23DB246DB6B6B6B6B5B6B66D2424641B9224B5B66D6D6D246D6D6D6D2423),
    .INIT_1A(256'hAD23D223FFFFFFFFFFFFFFFFFFFFFFFFFF6DD224DB9200D26C24DBDB24DB9224),
    .INIT_1B(256'h1BD2D2481B1BD289D2D2ADADD21B6C6423231B64ADACACAD646C6C6C646C6C6C),
    .INIT_1C(256'h25D31D1C1C65AE1CD41C1D6EAEAEF76E24F7FFFFDBD21BDA1BD264231B641B6C),
    .INIT_1D(256'hAE6EAEAE6565AEF7AEAEAE65AEAE6DAEAE6565651C6EB7AEAE6E6565AE1CD365),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFAEDC1C66AEAEAE6565656565656666652565666665656E),
    .INIT_1F(256'hFFF6F7FFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_006144_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i6_008,inst_doa_i6_007,inst_doa_i6_006,inst_doa_i6_005,inst_doa_i6_004,inst_doa_i6_003,inst_doa_i6_002,inst_doa_i6_001,inst_doa_i6_000}));
  // address_offset=7168;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFBFFFFFFFFFFBFEDFBFF2BF086EFFFFCFFFB3B39FFF3FFFFEFFFFFF),
    .INITP_01(256'hFFFFFFFFFF7FFFFFFFFFFDFF43FFF07F005C7FFFEFFFA7E67FEE7FFFFF7FFFFF),
    .INITP_02(256'hFFFFFFFFFEFFFFFF7FFFFEFFA3FFE46F0098EBFFE7FF4F9CFFDCFFFFFFBFFFFF),
    .INITP_03(256'hFFFFFFFFFCFFFFFF7FFFFF3F83FFE46E003197EFE7FF3E33FF39FFDFFFDFFFFF),
    .INIT_00(256'h6DAD6D246D6C24DB6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h24DBDB64B6B6B6B6B66DB6B664232424DB9224B5B66D6D6D6C6DAD24AD6D6D24),
    .INIT_02(256'hADACDA49B6FFFFFFFFFFFFFFFFFFFFFFF6DA231B9200246D24DB2424DB926DB5),
    .INIT_03(256'hD28989921BDA89D2D2236CD21B6C63DA1A1B64ADADADAD646CADAD64636C6CAD),
    .INIT_04(256'h251CD31C1C1C6E651CDC1C256EAEAEF76D24FFF648DA1BD21BDA641B1B236464),
    .INIT_05(256'hAEAE6E65AE6D65AEF7AEAEAE65AEAE65AEAE256565DC65AEAEAE6E6565AE1C8A),
    .INIT_06(256'hFFFFFFFFFFFFFFFF6D931D6EAFAEAE6D656565656565656665256566666E6565),
    .INIT_07(256'hFFF7F7F6F6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h64ADB56424AD6C24DB6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h9223ADB6B6B6B66D6DB66DDB232424DB926CADB6B66C6D6C64B56C24AD6D6D64),
    .INIT_0A(256'hADAD23401BFFFFFFFFFFFFFFFFFFFFFF24DB24DA926D6D2424241B92DB6D6DDB),
    .INIT_0B(256'h898989D2DB9191D2DA64D21B6C1BD2D2D264B5AD64642364ADAD6C631B6CADAD),
    .INIT_0C(256'h8B1CDCD3D4DC65AE65251C1C256EAEAEB76D652489DADADADA1B641B1B1B6423),
    .INIT_0D(256'h6EAEAEAE65AEAE65AEF7AE6EAEAEAE6565AEAE1D6566D41DAEAE66666565AE1C),
    .INIT_0E(256'hFFFFFFFFFFFFFF658A2566AEAEAEAE6D656565656666666E651D66656E65AE1C),
    .INIT_0F(256'hFFFFF6F6FFFFFFFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h646DB66D246DB56424DBB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h6CB6B6B6AD6D6CB5B624DA242424DB926D6DB5B6246D6D6C6DAD2323AD6D6D6D),
    .INIT_12(256'hACAD649149FFFFFFFFFFFFFFFFFFFFB6D224DBDB6D6D232424D292246D2492D2),
    .INIT_13(256'h499189D2D289D2D21BD2D2641B9289D264AD64DA1BDA23AD6C64641B1B6CADAD),
    .INIT_14(256'h1C931CD3D3D325656E65651C1C2566AEAEB66D92D21BDAD2DA1B64D21B23641B),
    .INIT_15(256'hDCAEB6B6AE65AEAE656DF7AE65AEAEAE6525AE651D6566D31CAE6E65651C65AE),
    .INIT_16(256'hFFFFFFFFFFFF25411C656EAE6DAEAE66666666666666666E651D6565AE65AE65),
    .INIT_17(256'hFFFFFFFFFFFFFFFFF6F7F7FFFFFFFFFFAEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h646DB5B6246CB66D6D24DBB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFEB66D6C246DB66DD2DA242424DBDA6D6DADB62464AD2464AD6DDB24B56D6D6D),
    .INIT_1A(256'h6CAC64D200B6FFFFFFFFFFFFFFFFFF24DBDB24B56C2424DB92DB2424DB921BB5),
    .INIT_1B(256'h898989D289D2D2D2D28923239291911B64D2D21BD21BAC64231B63D21BACADAC),
    .INIT_1C(256'h66D4D3D4D38B1C6D6E6565661C1C2565AEB66D89D21BD2DAD26423DA1B2364D2),
    .INIT_1D(256'hD324AEB6B7AE1CAEAE6565B7AE65AEF7AE1C1D66651D6566D4D4656665251C65),
    .INIT_1E(256'hFFFFFFFFFF6541D41DAEAE656EAEAEAE6E6E65AE656665AEAE1C65AE65AE65AE),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFF6F6F6FFFFFFFFB66DFFFFFFFFFFFFB6B6B6F7FFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_007168_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i7_008,inst_doa_i7_007,inst_doa_i7_006,inst_doa_i7_005,inst_doa_i7_004,inst_doa_i7_003,inst_doa_i7_002,inst_doa_i7_001,inst_doa_i7_000}));
  // address_offset=8192;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFF9FFFFFFBFFFFF9EC1FFE46E00212F6FE7FE7867FC73EFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFF3FFFFFFDFFFEFCFF0FFE0FE000078CFE7FEE19FF9E7DFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFE77FFFDFDFFFF6E770FFC0DC0000618EEFFDC33FE79FB7FFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFE4FFFFDF6FFFBB73B87FC0DC001B8A5DAFFF06778F3F6FFFFFFFFFFF),
    .INIT_00(256'h646C6DF66D24B6B66D6D2324FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hAD642464B56DDB92DB246424D2DB6D6DADF624DBB624656D6D641B64B56D6D6D),
    .INIT_02(256'h646464DB006DFFFFFFFFFFFFFFFFB6DBDB6DAE64249292D2DB241B92926DFFF6),
    .INIT_03(256'h9192899289D2D2D289D223D29289DA1B91D212D11B641B1BD2641BD21BADF564),
    .INIT_04(256'h6565DCD3D3938B656E6E6565651C1D2566B66489D21BD2DADA641BDA1B642489),
    .INIT_05(256'h658B65AFAEB7AE1C6E6E6565AEAE25AEF6AE1C1D655D1D6666D4D46565651DDC),
    .INIT_06(256'hFFFFFFFF6642D41CAE6D1CAEAEAEAEAEAE6666AE65AE65AEAE1C65AE65AE6565),
    .INIT_07(256'hFFFFFFFFFFFFFFF6F6F6AEFFFFFFFFB6FFFFFFFFFFADADAEB6B6F6FFFFFFFFFF),
    .INIT_08(256'h6D246DB6B6246DB6AD6D6D246CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h24246DB52491DA246C6D1C92DB6D6CB5F66492B66C24256D64631B64B66D6D6D),
    .INIT_0A(256'h646364DAD264FFFFFFFFFFFFFFFF24DB6DB624DA0000921B24DB911BB6FEAD24),
    .INIT_0B(256'hD292929289D292D289DBDA899192D291D21B1B5B1BDADA891B1BD1D223B5AD1B),
    .INIT_0C(256'h1C65251C93D38BD4666D6E2465661D1D25651B89DADAD2DB1B641A1A1B641B89),
    .INIT_0D(256'hAE1CD466AEAEF7AE1C6E666565AEAE1D6DF76ED41D1D1C1D6625D3D31D1D1D1C),
    .INIT_0E(256'hFFFFFFB641D41CAE651CAEAEAEAEAEAEAE65AE6E65AE656EAE1C65AEAE66AE1C),
    .INIT_0F(256'hFFFFFFFFFFFFF6F6F7F6F6FFFFFFFFB6FFFFF6FFFFB6B6FFFFFFFFFFB6FFFFFF),
    .INIT_10(256'h6D246DB6F66D24B6B66D6D6D24B5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h6D6D6C9292236C6D64DB92236424B5B624896DADDB246D6D63641B6CB56D6CAD),
    .INIT_12(256'h641B23922464FFFFFFFFFFFFFFB6926DB624DA0000921B2493922CB6B6641B24),
    .INIT_13(256'hD29192899191919291DA8989D2D289D1DA641BD289D1911B1BD291DA63B563DB),
    .INIT_14(256'hDC1C6565D4938B8B25AE6D656566AE25651C89D2DADAD2DB1B63D21B1B64DA89),
    .INIT_15(256'h65668B1CAEAEAEF7AE1C65656565AE661C65F765D41D25DC1D651C93D31C1D1C),
    .INIT_16(256'hFFFFFFD38B14651CD3AE6EAEAEAEAEAEAE65AE6565AE656EAE25DCB7AE65AE1C),
    .INIT_17(256'hFFFFFFFFFFFFF7F6F6F6F6F6FFB6B6F6FFFFFFB6B6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h6D246DB6F6B524ADB66D6DB66D24FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h6DDB49DB646D6D1BD2D2242424B6B523496DB6DB24246D2464641B6D6D6D646D),
    .INIT_1A(256'h1BD264D2246DFFFFFFFFFFFFFF246DB6DBDB9200D2241C92DB6DB66CDB1B646D),
    .INIT_1B(256'hDA91D28991919192D2D1891A12881AACADD100D21BD21AD2911BD21A64ACD21B),
    .INIT_1C(256'h1CD41C651D8B938BD465AE6E656566AE651C92D2DAD2D2DB241BD21B2364D2D2),
    .INIT_1D(256'hD366258A1CAEAEAEF7AE1C1C251D1C6666D465AF25D31C1DD425651CD3D31C1C),
    .INIT_1E(256'hFFFF2541D41CD3D3AE656E6E6EAEAEAEAE65AE656EAE656EAE658BAEF7AE6E6E),
    .INIT_1F(256'hFFFFFFFFFFFFFFF6F6F6F6FFFFF6F6FFFFFFFFAEB6AEB6B6B6FFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_008192_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i8_008,inst_doa_i8_007,inst_doa_i8_006,inst_doa_i8_005,inst_doa_i8_004,inst_doa_i8_003,inst_doa_i8_002,inst_doa_i8_001,inst_doa_i8_000}));
  // address_offset=9216;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFC9FFFFDFA7F7DDB1987F81DC0037BCDDAFFE48EF3C7CDFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFF93FFFFCFB3F8EE980C3F81DD003FFF99BFFED1BC707DDDFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFF83FFFFEFD9FC02080E3F8199007FFFA1BFF4A321E0FFAFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFF87FFFFEFC8FC8100071F819901FC1F037FFC44C7C3FF5BFFFFFFFFFF),
    .INIT_00(256'hB5246CB6F6B6646CF6AD6D6DB66D6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h92DB246D6D24DB92DB1B236CB56DDB9224B6DB23246D2C23A4A41B6D6D6D646D),
    .INIT_02(256'h1B926CDB6CB6FFFFFFFFFFFFB6246DDBDA23899224DB92DB6D6D23DB246D6C23),
    .INIT_03(256'hDA91D29191929192D2891264D11AEDF5ACDA6CADED5B88D1631BD21B641BD21B),
    .INIT_04(256'h1CD4D41D25D48B8B8A1C6DAE6565656EAEDB8AD2DAD2DA1B641BD21A646489DA),
    .INIT_05(256'h1DD365DC8B1DAEAEAEF7AE1CD31C1C1C2666D365AE1CD31C1C93651CD3CBD314),
    .INIT_06(256'hFFB641D41CD341AEAE65AE65AEAEAEAE6665AE1C6EAE656E65AE9325B7AE65AE),
    .INIT_07(256'hFFFFFFFFFFFFFFFFF7F6B6F6FFFFFFF6FFFFFFB6F7B6AEB6ADB6FFFFFFFFFFFF),
    .INIT_08(256'hB52424B6B6B66D24B6B66DADB6F624B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hDB246C24DBD2D2DBE4246C6D2423DB24B624DB24246CDB6CA49B1B6D6D6D646D),
    .INIT_0A(256'h2392AD23ADB6FFFFFFFFFFFF242424921B1BD224DB92DB2C24DB1B6424249292),
    .INIT_0B(256'hD291D29292D29191D28964A463F5F5F5ACF5F6F6A41A63F5ACD1D21B1BD2D223),
    .INIT_0C(256'hD4D4D3DC1D1DD48B4AD365AE6E6565656DD392D2DAD2DA1B641AD21B641B891B),
    .INIT_0D(256'h668B1C658BD31DAE6E6EAFAE1C8AD3D31D1D25D31C651CD31CD4D3651CD38BD3),
    .INIT_0E(256'hFFDC8A14D40165AE65AE6565AE66AEAE6565AE1CAEAE656E65AEDCD3AEF76E66),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFF7F7B6F6FFFFFFFFFFFFF6ADFFFFB6FFFFFFFFF6F6FFFFFF),
    .INIT_10(256'hB52424B6B6B6AD1BB5B66D6DADFFB56DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h6D641BDBDADADADB242C241B642324AD24DB24DB64231BEDA45B646D6D6C646D),
    .INIT_12(256'h1BD2F624FFFFFFFFFFFFFFB6DB64DBDB23DB24DA49DB2424DBDB1BDBDB92DB6D),
    .INIT_13(256'hD2D2D291D2D2D2D2D21AACEDECEDF5ADADB5F5F5ACF5F6F55B891BDB92D2D26C),
    .INIT_14(256'hD3D4D3D31C1C1DD38A421C65AE661D65248AD2DADAD2DA1B64D2D21B64DAD21B),
    .INIT_15(256'h6E1D41651D8AD41D666665AE6E1C93D3CAD3DCD44AD41C8B8AD342DC1C93938B),
    .INIT_16(256'hAE01D4D441D36E6566AE1D6EAE66AEAE1D6EAE1CAEAE65AE256E1D8A65AEB765),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6F6F7FFFFFFFFB6FFFFFFFFF6FFFFFF),
    .INIT_18(256'hB52423B6B6B6B51B6DB66D6DB5B6FF24B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h641BDBDBDBDB1B24641B1B6D24236D23DA24DB2464926CEDA35B642C6D64646D),
    .INIT_1A(256'h406DFF6DFFFFFFFFFFFFFF242424DBDBDB239A00DB24DBDB2424DBDBDB2C6D6D),
    .INIT_1B(256'hD2D2DA89DAD2DA1A5BA4F5F5F56489924991D264F5F5F5AC89D2D289D24824B6),
    .INIT_1C(256'h8BD4D38BD41C1D1D418A8A1D6EAE251C1B92D2DAD2D2DA2464D2D22364D2DA1B),
    .INIT_1D(256'h6565CB8B1DD48AD41D656565661CD38913D38AD3DC93D41D938BD342DCD48A8A),
    .INIT_1E(256'h1C8AD48A42656565AE6E1CAE656EAEAE1CAEAE1CAEAE1CAE1C66658A1CAEF7AE),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFB6FFB6F6B6B6F6FF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_009216_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i9_008,inst_doa_i9_007,inst_doa_i9_006,inst_doa_i9_005,inst_doa_i9_004,inst_doa_i9_003,inst_doa_i9_002,inst_doa_i9_001,inst_doa_i9_000}));
  // address_offset=10240;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFF07FF7FE7E47EED84030E139A03FE0F077FFC8BCF877E97FFFFFFFFFF),
    .INITP_01(256'hFFFFFFFE0FFF7FF3E22F7804038713BA0BFE0FAFFFF8D7FF9DFDB7FBFFFFFFFF),
    .INITP_02(256'hFFFFFFFE3FBF7FB3E0013C0001C703320BFE3F7FFFF3CDFF87FF7FFBBF7FFFFF),
    .INITP_03(256'hFFFFFFFE6FBF77B1F0003E0001C303360BFE3FFFFFF387FE1F3FFFFFBF7FFFFF),
    .INIT_00(256'hB6241BB6B6B5B6236CB6AD646DB6FFB66DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h1BDADBDBDB24241BD264AD24246D23DA24DBDB24DA23F5ECA35B6D246D246464),
    .INIT_02(256'hDBFFF6F6FFFFFFFFFFFFB6236C1BDBDB1BD200DB24DB2364231BDBDB6D6D641B),
    .INIT_03(256'hD2D2DA91DBD21A63ACECF5EC5B231B00000000006CF6F51B889289D24023F624),
    .INIT_04(256'h8B93D38BD3D41C6593424AD365AEAEDB92D2D21BD2D21B641B91D26464911BDA),
    .INIT_05(256'h65651C42D31D938BD41C1C1C1C1D1DD313A45BD2131CD41D1C8BD38AD31D8B8B),
    .INIT_06(256'h42D49342DC652565AE251CAE656EAE66DCAEAE1C65AE1CAE1D2566D38A65AEAF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6B6F6FFFFFFB6B6F6F6B6F6F76D),
    .INIT_08(256'hAD1B1BB6B6B5B62424B6AD6D64B6FFFF24B6FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h1BDBDB1B1B1BD21BADF5231B2424DB231BDB231BDBADF6A45B636C246DDB246C),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFF6D2424DBDBDB646C9224DB24241B1B1B646D641B6463),
    .INIT_0B(256'hD2DADA911BD21AA4F5F5F5F5B5FE6D004A4A49DA23FEAD1A1BDA1B9264FFB523),
    .INIT_0C(256'hD38BD3D38BD31C651C8A8A8AD465AE6589D2D21B89DA1B641B891A6C1BD223D2),
    .INIT_0D(256'hAE651DD341D41C8B8AD31CDC1C1D1D1CCA1BA4A312D3D4CBD4D38A8B4114D48A),
    .INIT_0E(256'h8BD38BD31D651C656E1C65AE6566AE65D3AE6E1C65AE1C66251C6E1C8ADC66AE),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6FFFFFFF6FFFFF7AEB6F6FFFFF7D3),
    .INIT_10(256'h6DDB23B66DB5B664DBB66D6D24B5B6FF6D6DFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h1BDBDBDBD21AA4F6B51B1B2364641B1BDB1B232323F6F5A35B64246C6DDB246C),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFB6246CDBDB1B64AC64DBDB2424DB232364641B5BAD641B),
    .INIT_13(256'hD2DADA921BD21AACF5F4F5F5F6FFB6DC4A0024FEFEFEF5ADDA241B6DFFFFB5FF),
    .INIT_14(256'h8B8B8BD3D3D3D465651C8A8A8A1CAE6592D2D2DA91DA1B64D2891B6CDADA1B89),
    .INIT_15(256'hAE6E25D48A42D4D48A8AD3D4D3D3D41DD4D25BA3A35BD2D38BD4D38A8A8ADC8B),
    .INIT_16(256'hCB8B1C1C651D1D6E6ED365651D65AE25D3AE661C1CAE1C6565D365258B8B2565),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFF6FFFFB6B6F6FFFFAE8A),
    .INIT_18(256'h6DDA24F66DB5B664DBB66D6D246DB6FFFF6DFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hDBDBDB1B64F5F6ACDBDB24AD6C1B1B1B1B1B642364F5A3635B641B6D2323246D),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFF652424DBDA24B51BD2DBDBDB1B2323232364ACA4641BDB),
    .INIT_1B(256'hDADAD2D21BD21BACF5F5F5F5FEFF259B49DCF6FEFEFEF66C236464F6FFFFFFFF),
    .INIT_1C(256'h8AD38BD3DCD3D3256525D3D34AD3651CD2D2DBD2D2DA236492896464D21B1B92),
    .INIT_1D(256'h656E661DD38A8AD3D38B8AD3D4D3D3D4D4D31BACA3A35BD28A8BD38A8A42D3D3),
    .INIT_1E(256'h8B1C65DC1D1C1D6E669365651D65AE1CD3AE651CD4AE1C1C65D31C65D38BD365),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAE41),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_010240_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i10_008,inst_doa_i10_007,inst_doa_i10_006,inst_doa_i10_005,inst_doa_i10_004,inst_doa_i10_003,inst_doa_i10_002,inst_doa_i10_001,inst_doa_i10_000}));
  // address_offset=11264;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFE6FBF7698F0001F8009C023350BFF7FFFFFE305F83EFFFFF7BF7FFFFF),
    .INITP_01(256'hFFFFFFFCDFBF62C8FB300F8009C007754BFFFFFFFFEEE3C03BEFFFB7BF7BFFFF),
    .INITP_02(256'hFFFFFFFCDFBE6A48791800000CE0066D4BFFFFFFFFCDE7800FFFFFB73F7BFFFF),
    .INITP_03(256'hFFFFFFFCC3A668041D9C00000DE0466B4BFFFFFFFFD9EF803FFFFF7B3F7FFFFF),
    .INIT_00(256'h64D224B66DB6B564DBB56D6C2423B6FFFF6DB6FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h4A9264B5FEF523D2236DF6AD1A1B241B1B646C23F5AC5A1A1B24236DDB24236D),
    .INIT_02(256'hFFFFFFFFFFFFFFFFB6246DDBDADB6C6CD2DBDBDBDB24DB2364AC646C23DBDBD2),
    .INIT_03(256'hDBDBD2D21BD25BACF5F5F5F5FE6C1C24DBF6FEFEFEF6636423646CB6FFFFFFFF),
    .INIT_04(256'h8A8B8B8B1CD3D31D6665D4D38B4ADBD3D2D21B92D2DA646489D26463D223D21B),
    .INIT_05(256'h25656665D4D2D38AD4D4D381CBD4D3CBD3D48AA5F5A3A363138AD3938A4A8BD3),
    .INIT_06(256'h8A6E65D41C1C1D66658B651D1C65661CD3AE651CD3651DD465DC8B651C8A8BDC),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFFFFFFFFFFFF1C42),
    .INIT_08(256'h24926DB624B6B564D2ADAD246CDBADFFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h01001AB56CDA236DF6FEADD21B6C231AACAD23ADF6ECAC631BDB2464DB2423AD),
    .INIT_0A(256'hFFFFFFFFFFFFFFFF6D2424921B641BD21A2423DBDBDB2363ED64409293924949),
    .INIT_0B(256'hD21BD2D21BD263ACF5F5F5F6FE1B1B24ADFEFEFEF663646C1B6464F6FFFFFFFF),
    .INIT_0C(256'h8B8B938A1DD48B1C6565D48BD48A8AD2D2D2DB89D21B641B401BAD1BD263D21B),
    .INIT_0D(256'h1C1C65661D8A1B138AD31C1B898BD3D3CBD3D3D3ADED635B5CD38AD38B8A8AD3),
    .INIT_0E(256'h24F7D41C1C1C1D661D93651C1D1D651CD36665D4D4DC25D31D1C8ADC1D938A93),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFD342),
    .INIT_10(256'hDBD26DB524B6AD24926DAD246DDB6CB6FFFE6DFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h00DB92D264B5FEFEFEF51A64B56C1AADF56C64FEF5ACEC641BDB241BDB1B246D),
    .INIT_12(256'hFFFFFFFFFFFFFFB6246DDB9264249123A46424D2DB2424641B89004A49494A4A),
    .INIT_13(256'hD21BD2DA1BD263ECF5F5F6F6FEFE6D6DFEFEFEFE6463AD641BAC64B6FFFFFFFF),
    .INIT_14(256'h8B8AD38A1D1D8BDC65651C42D4D38AD3D2DADB89DA1B6CDA00646CDA1B1BDA1B),
    .INIT_15(256'h931C1C6665D3D25CD38AD36464898A8B8B8BD39392D29240898A418A934A8A8B),
    .INIT_16(256'hB6B642141C1C1C661C93651C1C1D65DBD36565D31CD31CD3D41D938B1CD48A8B),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAE8A42),
    .INIT_18(256'hDADBB6646DB66D24D26DAD246D2324B6FFFF6DFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h00DB6DB6FEFEFEFEF5636CF6AD1AB5F6AD23FEFEEDECF523DB246C1B1BDB6464),
    .INIT_1A(256'hFFFFFFFFFFFFFF6C642492246CDAD2B5E46323D21B24646D6D49008A8A8A4A52),
    .INIT_1B(256'hDA1BD2DA1BDA63F5F5F5F6F6FEFEFEFEFEFEFEF66C6C6D241BAC64FFFFFFFFFF),
    .INIT_1C(256'h8B8A938A1D258B1C656E1D4AD3D3D3D3D21BD292DB2364D1886C64D223D21B1B),
    .INIT_1D(256'hD38BD41C651C8A1B64CA4113AD63D28B8B8B8B8B8A00000000000041934A4A8A),
    .INIT_1E(256'hFF658BD4D4D41C661C8B25DCD41D65D3D36565D31C8BD4D38BDCD48BD31C8BD3),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6D41D4),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_011264_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i11_008,inst_doa_i11_007,inst_doa_i11_006,inst_doa_i11_005,inst_doa_i11_004,inst_doa_i11_003,inst_doa_i11_002,inst_doa_i11_001,inst_doa_i11_000}));
  // address_offset=12288;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFDC3A660008CCF00000DE0466ADBFFFFFFFF99EFE07FFFFFF37F7DFFFF),
    .INITP_01(256'hFFFFFFFD83226040C66600000DE04EF2DFFFFFFFFFB3EFE07FFFFFF67E7DFFFF),
    .INITP_02(256'hFFFFFFF983332040637980000DE09CD45FFFFFFFFF73EFE27FFFFFE67E7DFFFF),
    .INITP_03(256'hFFFFFFFB83333060713D80000DF09CC45FFFFFFFFF66CF93FFFFC3E4DDFDFFFF),
    .INIT_00(256'h9224B523B5B66424DB6CAD246D6CDBB6FFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h0024FEFEFEFEFEF6ADB5FEB51BB5FEF664F5FEF6F5F66C1B1B246464DADB6D1B),
    .INIT_02(256'hFFFFFFFFFFFFB6246DDBDB6D2392DAADAD2324DA232464ADF5ADB6DC498A4A8A),
    .INIT_03(256'h1A1BD21B1BDA64F5F5F5F6FEFEF6FEFEFEFEFEF6F5ACAD241B6C64FEFFFFFFFF),
    .INIT_04(256'h8B8A8B8A1C65D31C6566658B8BD3D2D2D21B89D2DB646440D26D23DA239223D2),
    .INIT_05(256'h5BCA8BD31C65D4CA5BA3D2011CEDAC1A014A8B8B8B8A4941828242018A8A4A8B),
    .INIT_06(256'hFF1C93D4D4D41C651C8B25DCD41C65D48A1D65D3D4938BD3D2D3D48B8BD3D3CB),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF25006D),
    .INIT_08(256'hDB6C6C23B6AD24DBDB64AD246D6DDB6DFFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h00ADFEFEFEFEFEF6F6FEB523F6FEFEACADFEF6EDF5F523642424AD23DB2424DA),
    .INIT_0A(256'hFFFFFFFFFFFF246D2492246D92DA1B6CAD2423DA242464ADADF6B69B4A8B8B8A),
    .INIT_0B(256'h1A1BD21B1B1B64F5F5F5F6FEFEFEFEFEFEFEF6F5F5AD64641B6C64FFFFFFFFFF),
    .INIT_0C(256'h8B8A8B8A1D65D31C1D6E65D38A8BD2D2D21B89DB1B6C230023AD1B1BDADA1BD2),
    .INIT_0D(256'h1B5C8A8BD31D1DD3D2A4A4D20064ED88018A4A8B8B8A414141414141418A8A8A),
    .INIT_0E(256'hFFD3D3D3D4D31C65D48B1DDCD3D41DD48A1C65D38A8B8BD3D313D3D38A8AD38B),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1C00FF),
    .INIT_10(256'hDB6D1B64B66D1BDBDB246D2464B6DB6DFFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h00F6FFFEFEFEFEFEFEF66CF6FEFEB5ACFEF56C64AC63646C1B64B5DBDB241BD2),
    .INIT_12(256'hFFFFFFFFFFB6246DDA246D2392DB24646C641BDB24246CADAD646EDC010225DC),
    .INIT_13(256'hDA1BD21B1B1B64F5F5F6FEFEFEFEFEFEFEFEFEF6F6AD641B1BAC64FFFFFFFFFF),
    .INIT_14(256'h8A8A8B8A1D66D41C1D6566D441D3D3D11BDA911B1B6CDA00646CDA1BD21BD2D2),
    .INIT_15(256'hD2A45C8A8BD31C148A1BA4A41B41D2636E9201418A8B424141414141004A8A8A),
    .INIT_16(256'hF792D3D4D3D31C65D48B1C1C8BD41D1C8BD465D38AD38B93D31BD3D38A8A8AD3),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF93DBFF),
    .INIT_18(256'h2424DBADB624DB1B23246D2424FEDB24FFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h24FFFEFEFEFEFEFEFEF6FEFEFEF5ACFEF61B490092DB6C231BF66C92DC24DADB),
    .INIT_1A(256'hFFFFFFFFFF646D1BDB6D6D92D22364DB2464DBDB24246CADAD00DC6F01936E2D),
    .INIT_1B(256'hDA1BD21B1B1B64F5F5F5FEFEFEFEFEFEFEFEFEF6ACAC6C1B1BAC64FFFFFFFFFF),
    .INIT_1C(256'h8A8A8B8A1C66DC1C1C65661C41D3DBD11BD2D21B636C8992AD64DADAD21BD2DA),
    .INIT_1D(256'h8B1BAD5BCA8AD31CD4CA63A3EC650064B6920041938A8A4141414141004A8ACB),
    .INIT_1E(256'hF78ADCDC8BD31C1DD48A1C1C8BD31C1C8B8B1C1C4AD3D38A8A1C1CCA8AD48ACA),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF006EFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_012288_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i12_008,inst_doa_i12_007,inst_doa_i12_006,inst_doa_i12_005,inst_doa_i12_004,inst_doa_i12_003,inst_doa_i12_002,inst_doa_i12_001,inst_doa_i12_000}));
  // address_offset=13312;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFBB11132323C1ED80007F09DC8DFFFFFFFFEE6CFBCFFFF01C8B9FDFFFF),
    .INITP_01(256'hFFFFFFFBB11013333E1FB80407F9BDCAFFFFEFFFFCCCCFC0FFFF00C1B9EFFFFF),
    .INITP_02(256'hFFFFFFFFB000113B9F8FF84607F13986FFFF9FFFFDCCDFF7FFFFC00371EFFFFF),
    .INITP_03(256'hFFFFFFFFB000018DEFE7D86607F17B86FFFFDFFFFB9CDFFFFFFF810071EFFFFF),
    .INIT_00(256'h24DB24B66DDBD21B24246D2324FFDB24FFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hF6FFFEFEFEFEFEFEFEFEFEFEFEF5FEFEDB004A4A4A00DA1BACF5DBDB24DBDADB),
    .INIT_02(256'hFFFFFFFFB66464DA246D2492DB6424D21B64DBDB246CADADF6D225B76E6EDCDB),
    .INIT_03(256'h1A1BDA1B1B1B64F5F5F5F6FEFEFEFEFEFEFEFE6463AD641B1B6C64FFFFFFFFFF),
    .INIT_04(256'h8A8A8B42DC6E1C1C1C66662593D3D2DA1B89DB1B6464001BAD1BDA921BDAD2D2),
    .INIT_05(256'h8BD3A4ECA4138A8BD48BD2A4ECEDADD26C1B41F765008A824182824200DB93CB),
    .INIT_06(256'hF78A1C1C8BD3D41CD48BD41C8BCBD41C934A1C1D428A1BD34AD3641281D41C81),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF701B7FF),
    .INIT_08(256'h23DB6DAD24DA922464246DDB64FF2423FFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hF6FFFEFEFEFEFEFEFEFEFEFEFEFEFEF692924A4A4A4A9340AD64D2DBDBDBDB23),
    .INIT_0A(256'hFFFFFFFF246DDBDB6D6DDBDA246CDBDB1B6DD2DB246CADADF51B928ADC930092),
    .INIT_0B(256'h1B1B1B231B236CF5F5F5F6FEFEFEFEFEF6F66391ACAC641B1BAC64FFFFFFFFFF),
    .INIT_0C(256'h8B8B8B8AD3651C1C1C656E651BDBD21B1B911B236C1B00646C1AD2921BD21BD2),
    .INIT_0D(256'h81421CEDECA45CCA41D38A1BACECF5F56CDB6DFF25418B8282828A8A0024D3CB),
    .INIT_0E(256'hF74A241C4A8BD41CD48BD31C8BD3D3D4D38AD31C8B41131B428A5BA4D282651B),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6D3FFFF),
    .INIT_10(256'hDB1B6D6CDB92D2246D6D6DDB6DFF2424FFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hF6FEFEFEFEFEFEFEF6F6FEFEFEFEFEB6B625019349924A0092DBDBDBDBDB1B1B),
    .INIT_12(256'hFFFFFFAD6D24DB64B624DADB6C24DBDB246DD21B246CADADAC631B1BDB24646C),
    .INIT_13(256'h1B1B1B231B6364EDF5F5F6FEFEFEFEF664DA401AAC64641B1BAC64FFFFFFFFFF),
    .INIT_14(256'hD3D38AD3D3651D1C1C656E65D3DBD21BD2D22364ACD192AD64D291DADA1A1BDA),
    .INIT_15(256'h1A8A0165F6ECECED1B414A8A64ACACFEFE2465B76582CB828A1C8A41006D1C8A),
    .INIT_16(256'hF74A6565418BD4D4D4D38BD4D38B8BD3D48A8A1CCB8AD264D341136464CA13AC),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB624FFFF),
    .INIT_18(256'hDB646D1BDBDBDB6DB66D24DBADFF2424FFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFEFEFEFEFEF5F5F5FEFEFEFEFE6DB6DC414A4A4A0025DB92DBD2DBDBDBDB),
    .INIT_1A(256'hFFFFFE6D6DDB23B56DDBDB246D23DBDA246D92236C6CADEDEDF5F6F6FEFFFFFF),
    .INIT_1B(256'h1B1B2364236364ACF5F5F6FEF6FEFEAC1A1A8923AD64641B1BAD64FFFFFFFFFF),
    .INIT_1C(256'hD4D38ADCD365651C1C656E6DD2D2DA1BD21B236464401BAD1BD291DAD21B1BD2),
    .INIT_1D(256'hEC641300ADF6ECF5F6AD13410064F5F5FEF74965F78B42D300AEAD0000B62541),
    .INIT_1E(256'hF74A6D6E41D3D3D4D4D38AD3D38B8BD3D4D38AD3D38AD2646441CAD21B1B89A4),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB66DFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_013312_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i13_008,inst_doa_i13_007,inst_doa_i13_006,inst_doa_i13_005,inst_doa_i13_004,inst_doa_i13_003,inst_doa_i13_002,inst_doa_i13_001,inst_doa_i13_000}));
  // address_offset=14336;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFB4000180F7FBECF697F37B0CFFFEDEFFFB98DFFFFFFE8308FDEFFFFF),
    .INITP_01(256'hFFFFFFFFF4000000FFFFE7FE97F2F31CFEFD9EFFF738DFFFFFFFB3C1BFFFFFFF),
    .INITP_02(256'hFFFFFFFFFE000000FFFFEFCE97E6F739FE71BEFFFF38DFFFFFFEFF82FBDFFFFF),
    .INITP_03(256'hFFFFFFFFDE000000FFFFE00E97E6F631FE01BEFFEE74DFFFFFFF1F25FBDFFFFF),
    .INIT_00(256'h24241B242424DBADB6AD24DBF6FF246DFFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFEFEFEFEFEFEF5F5ADADFEFEFEB6922D004A93920024B6DADBDBDB1BDBDBDB),
    .INIT_02(256'hFFFF6D6D24DB6DB524DBDB6D6DDBDBD2246DD21B6D6DADEDF5F5F5FEFEFEFEFE),
    .INIT_03(256'h1B1B64641B646464F5F5F6FEFEF663D21B1A89646C2364D223AC64FFFFFFFFFF),
    .INIT_04(256'h1CD38B1DD365651C1C656E65DBD21B1BD223636C23486C6CDA89D2D21B1BD2D1),
    .INIT_05(256'hEDECED6441ADFEF5F5FEF6AD1B896CF5F6FF6492ADAED3001BEEF71C49FF6541),
    .INIT_06(256'hFF926DB68A1CD393D3D38A8BD38B8B8B93D38B8BD38AD21B1C498A41009149DA),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6FFFF),
    .INIT_08(256'h24DBB5246D2424B6FFAD1B23FFFF246DFFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFEFEFEFEFEFEFEF5F5EDF6FFFEFE231C77DD256E00DBF7242423D2DBDBDADB24),
    .INIT_0A(256'hFFB66D6CDB64B66CDBDB246D24DBDB922C6DDB236D6DB5ADF5F4F5F5F5F6FEF6),
    .INIT_0B(256'h1B1B646C236464D2ACF5FEFEF51B891B1BD2D26C642464D264AC64FFFFFFFFFF),
    .INIT_0C(256'h1CD48B1DD325661C1C65651CDAD223D21B23646CD2D2AD64D292D21B231B91D2),
    .INIT_0D(256'h64F5F5F6AD24ADFEF5F6FEFEF6B664B5F6FFB600D3FFF765F7A55D6524FF6582),
    .INIT_0E(256'hFF1C65F7D325D48B8B938B8AD38B8B8A8B8B8B8A938A894100004A8A49000000),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6FFFF),
    .INIT_10(256'h1BF6B56DB6DB6DFEFF6DDB6DFFFF24B6FFFFB6FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hF6FEFEFEFEFEFEFEFEFEFFFEFEF62489256E261C1BFF6D6D6CDADADBDBDB1BDB),
    .INIT_12(256'hFF6D6D1B1BB5B524DBDB6D6D1BDBDBDA6C6DDB1B6D6DB5EDECF5F5F5F6F6FEFE),
    .INIT_13(256'h1B1B646C23646C89D1ACF5ACD248D21B1BD21B6C1B6464D364AC23B6FFFFFFFF),
    .INIT_14(256'h1DD48B1DD31D661C1C6565DBD21B1BD21B6364648964AC1B91921B641B92921B),
    .INIT_15(256'h1BF5F6F6FEF6ADF5FEFEFEFEFEFEFEF6F6FFFF921CEFAFEFA6134100B6FF648A),
    .INIT_16(256'hFF251CFF1C6525428B8BD38A8BD38B8A8B8B8B8A8AD289004141414A4A4A0100),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6FFFFFF),
    .INIT_18(256'hB6B624FFB6DBB6FFFF6D92B6FFFF24FFFFFFB6FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEF6F66D4900496DFFF6B6ADD2DA23DBDB1BDB24),
    .INIT_1A(256'hB56D24DB6DB66DDBDB246D64DB1BDBDA6D6DDB1B6DADADF5ECF5F5F5F6FEFEFE),
    .INIT_1B(256'h1B23646C2464ADD189D1898989D2D2231B8964641B6C1CD364AD232465B6FFFF),
    .INIT_1C(256'h1DD4D31DD31D661C1C6524DAD2231BDA23646423896C64D289DA6464D289DB1B),
    .INIT_1D(256'hADF6F6FEF5FEFEFEFEFEFEFEFEFEFEFEFEFEB68941CB418A404000926DB66D8A),
    .INIT_1E(256'hFFB6D3FF6D1CB68A8A8BD38A8A8BD38A8A8B8B8ACAD38A41414141428242418A),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_014336_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i14_008,inst_doa_i14_007,inst_doa_i14_006,inst_doa_i14_005,inst_doa_i14_004,inst_doa_i14_003,inst_doa_i14_002,inst_doa_i14_001,inst_doa_i14_000}));
  // address_offset=15360;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFDB000600FFFFF80697EDE663FE03BCFFDE78CFFFFFFFDE43FFDFFFFF),
    .INITP_01(256'hFFFFFFFFFF000230FFFFFFFE97EDECC27E036CFFFDF8CFFFFFFFFC8FFFBFFFFF),
    .INITP_02(256'hFFFFFFFFFF8003317FFFFFFE96EBEDD6FF0378FFBAFAEFFFFFFFFEBEFFBFFFFF),
    .INITP_03(256'hFFFFFFFFFFC001B9FFFFFFFE961BC9B6FF0658FF7FF4EFFFFFFFFDFFFFFFFFFF),
    .INIT_00(256'h6D24FFFF236DFFFFFF24DBFFFFFF6DFFFFFFB6FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEF62489B5FFFFAD92DB6CDBDBDBDB64B6),
    .INIT_02(256'hAD6CDB24B6B623DBDB6D6D2423DBDBDA6D6DDBDB6DB5ADACF5ECF5F5F6FEFEFE),
    .INIT_03(256'h1A646C6C6464ADD289898991D2911A641B92641B6464D3D264AC1B656524656E),
    .INIT_04(256'h1DD4D31DD31C661C1C251CD21A23D21B636464D2DA6C1B89926464D289D2231B),
    .INIT_05(256'hADFFFEFEFEFEFEFEFEFEFEFEFEFEFEF6F6FEAD641BD2D292D2D292D249ADAD8A),
    .INIT_06(256'hFFFF93FFFFD3F765018A8B8B428A938B8A8B8A8A8A1C1C004141418282824101),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h24F6FFB624B6FFFFFFDA6DFFFFFFB6FFFFB6FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFEFEFEFEFEF6F6FEFEFEFEFEFEFEFEFEFEFEAD6CFEB5DB9223DB92DB1C24B56D),
    .INIT_0A(256'hAD1B1BADB66CDB1B24AD6D2324DBDBDA6D6DDBDB6CB5AD63ECF5F5F5F6F6FEFE),
    .INIT_0B(256'hDA646C6D6464ADD2899192D2D2922364911B24DA641BD29264AC1C65656D2424),
    .INIT_0C(256'h1DD4D41DD31C661C1C1C1BD21B1BDA23636C64916364D289646CDB91D2DA64DB),
    .INIT_0D(256'h1CFFFEFEFEFFFFFEFEFEFEFEFEFEFEFEF6F5F5F6F5F5F5FDF6F6F6F6F6F6AD92),
    .INIT_0E(256'hFFFF24B7FF24AEFFD3418BD38A4A8A938A8A8A8A4A8B64D30000651D4142D341),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h24FFFF6D6DFFFFFFB6DBFFFFFFFFFFFFFFB6FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFEFEFEFEFEF5B5F5F6FEFEFEFEFEF6F6FEFEFEFEF6B61BD21BDB242324646DDB),
    .INIT_12(256'h24DB6DB6B6DB23DB6CAD24241BDB1BDA6DB51BDB6CB5B56363ECECF5F5F6FEFE),
    .INIT_13(256'h1A646CAD6423AD1B89D2D2D289DB641B491B1B2364DB92D264AC1B1C656525AE),
    .INIT_14(256'h1DD4D41D931C66D41C1B1BD264D2232364641BD1641B481BAD23891BDB1B24D2),
    .INIT_15(256'hD3F6FEFEFFFFFFFEFEFEFEFEFEFEF6FEF6F5F5F5F5FDFDFDFEFEFEFEFFFEAE92),
    .INIT_16(256'hFFFF6EAEFFF624FFF74141D38A4A8A8B8A8AD38A8A4113659200F7AE4141D3A5),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h24B6B624FFFFFFFF6D6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFEFEFEFEFEFEF6F6FEFEFEFEFEFEFEFEFEF6FEFFFFAD89246D24241B1B246D6D),
    .INIT_1A(256'hDB24B6B6241B23246D6D2424DB23DB926DB61BD264B6ADACA3A3F4F5F5F5F6FE),
    .INIT_1B(256'h1A646CAD6C1BAD6489DAD289D26C6489D21BD26423D28A9264AC1B1C1D1C6E6D),
    .INIT_1C(256'h1DD4D41D931C66D4D4DBD21B64D264236C64DBDA6489D2AD64896464D2641B92),
    .INIT_1D(256'h1CADF6FEFFFFFFFFFEFEFEFEFEFEFEF5FEFDFDFEF6F6F6F6FEFEFEFFFFFFB692),
    .INIT_1E(256'hFFFFFF6DFFFF6DB6FFB74241D38A8A8BD38AD3938A8A405CAD9224AE1C41D3EE),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_015360_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i15_008,inst_doa_i15_007,inst_doa_i15_006,inst_doa_i15_005,inst_doa_i15_004,inst_doa_i15_003,inst_doa_i15_002,inst_doa_i15_001,inst_doa_i15_000}));
  // address_offset=16384;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFE000CF7FFFFFFE96DFDB6CFB0CB8E6F5F4EFFFFFFFF9EFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFF800767FFFFFFE96B7D6EDFF1878E6EFFCEFFFFFFFFBDFBFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFC0170FFFFFFFE96B7DDD9FFB076EDEBECE7FFFFFFF79DFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFE027BFFFFFFFEB66F9DD3FFE0F2DBDFFCE7FFFFFFF7BDFFFFFFFF),
    .INIT_00(256'h6D6D6DFFFFFFFFFF24FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFDBDAB56C241BDB246DB6B6),
    .INIT_02(256'h246DF66DDB24DB6C6D6D2424DB24DB926DB623D223B6ADA4E49BACF5F5F5F6FE),
    .INIT_03(256'h64646CAD6CDAADADD1D28989646CD2891BD2236423928A9264AC1BD3D324ADDB),
    .INIT_04(256'h1DD4D41D931C65D31B1BD2641A1B6423AD64D21C1B89AC6C9225B6DB1B64D2D2),
    .INIT_05(256'h0024ADF6FFFFFFFFFEFEFEFEFEFEFEFEFEFEFEF6F6F6F6FEFEFEFFFFFFFFB6D2),
    .INIT_06(256'hFFFFFF6DFFFFFF6DFFFFB79200928B8B8B8B8A8B8B8B8B4164AD924A65AEEE65),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hB6DBB6FFFFFFFFB66DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFF6C916DAD2424DB1B6DB624B5),
    .INIT_0A(256'h6DB6B6DB2424236D6D2424232424DB9264B623DA1BB5B5ACECE39AECF5F5F5FE),
    .INIT_0B(256'hFF6D64ADB52463ADD20089646CD289D2DA1B64641B928A8A646C1BD3DBAE24DB),
    .INIT_0C(256'h1DD3D41D8B1C65D31BDB1B64D16423646C1BD21BD2646C9224B665D2641B8964),
    .INIT_0D(256'h0064ADACFEFEFFFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFB692),
    .INIT_0E(256'hFFFFFFB6B6FFFFB7B6FFFFFF1C00428B8A8B8A8AD38BD4D34064F61341AE6500),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hB624B6FFFFFFFFB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFB5D21BB66D6CDBDB24AD6D926D),
    .INIT_12(256'hB6F664DB64DB64AD6D2364DB6424DB9264B624DAD2B5B5ACECE3E39AECF5F5FE),
    .INIT_13(256'hFFF664ACADAD1BAD6489AD64D2D2D2DAD2232364D21B1C9223641B8A6D6DDB24),
    .INIT_14(256'h1DD3D41D931D65D31BD2641BD2641B6C641BD21A1B6CD21C6E6EDB1C64D2DAF6),
    .INIT_15(256'hACF6F5ACF5FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFB68A),
    .INIT_16(256'hFFFFFFFFFFFFFFFFB7FFFFFFFF6E8A428A8B938A8A93DC1CCA12ACEDD2410092),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hB66D6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFF6D23DB6DB56D24DB236DB56D496D),
    .INIT_1A(256'hF66DDB64241B6D6D242464236D24DB9224B62492496DB5ACECEBE3A39BEDF5F5),
    .INIT_1B(256'hFFFFAD64ADB564646D1C6491D2DAD2D21B1B6C23D2D31CD22464DB64AEDB246D),
    .INIT_1C(256'h1DD31C1D8B2565D2D21B64D223641BAD24D2D21A641BD365AE24D224D2926DF7),
    .INIT_1D(256'hFEFEF5F5FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFAE8A),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF6E008A8AD4D38A8B1CD4005BACED5B0064F5),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_016384_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n28 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i16_008,inst_doa_i16_007,inst_doa_i16_006,inst_doa_i16_005,inst_doa_i16_004,inst_doa_i16_003,inst_doa_i16_002,inst_doa_i16_001,inst_doa_i16_000}));
  // address_offset=17408;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFE01FFFFFFFFFEB66F9BB7FFC1E0FFF7FCE7FFFFFFDF3DFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFE07FFFFFFFFFEB6DB136FFFC3DCFFB7F867FFFFFE0F7DFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFE1FFFFFFFFFFEB6DB16ED8FE7FE6F6FF8637FFFF85E7CFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFE3FFFFFFFFFFEB7FF1DBFF7F7BEDFCFF8633FFFC73CFCFFFFFFFF),
    .INIT_00(256'hF6B624B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEF6AD23DB1B24B66D6DDBDB246DB66D9224),
    .INIT_02(256'hB6242464DB246D6D246C24246D23DBDA23B665920065B6ACECECEBEBA39BEDF6),
    .INIT_03(256'hFFFFF66C6CB5AC246D1C4ADBDBD2911B1B6464D2DB8A8A8A236423AE1C246CB6),
    .INIT_04(256'h1D8B1C1D8A6565D3D2642392641B23AD1B91D21B6492256E65D21B1BDBADF7F7),
    .INIT_05(256'hF6F6F5FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFAE8A),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFB74A8A8AD4D4D48AD31C6564ECF4ACADF6FE),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hB6FE24B5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEB564DB92DBDBDBADAD6D24DB236D6DB6AD9224),
    .INIT_0A(256'h64DB6C1BDB6D6D6D246D236D6CDBDBDADBB665920024B664ACECECE3E3A39BEC),
    .INIT_0B(256'hAEAEADAD6C6CAD646C244ADCDB891B231BADDB1B1B1BD38A2423AD241B24B6B6),
    .INIT_0C(256'h1C8B1C1C8B6565D21B6CD21B64D26C6CDA91D21BDBDB6D65D31B1BD264ADADAE),
    .INIT_0D(256'hF6F6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFFF6D8A),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7D38B8BD48B931C6EB7FFADACECF4F5F5F5),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hB5FF6D24FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hACF6FEFEFEFEFEFEFEFEB66C23DBDBDBDB23D26CB6AD6DDBDB246D6D6DB692DB),
    .INIT_12(256'hDB2464D21B6D6D24246D246D24DBDBDBDBB56D9201DBB624D2A4ECECEBEBA35A),
    .INIT_13(256'h13D3CAD36CACACAD64642449491B631BAD231B241C6565D3D26D6DDB24B5F66D),
    .INIT_14(256'h1D8B1D1C8A65658A6464D26464D2AD64D291D21BDB2465DB1B5B12CA1313D213),
    .INIT_15(256'hF6F6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFFF6D8A),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7D38B93D31CAEB7B7FFFFB664F4ECF5F5F5),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h6DFFB624B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hA3A4F5FEFEFEFEB56C23D292DB231B1BDBDB23B5B66DDBD22364AD246DB5D2DB),
    .INIT_1A(256'h1B6DDBD2246D6D236D64246D24DBDBDBDB6D6D8A024A6E6D004A1B64ACECECAC),
    .INIT_1B(256'h5CA5A513CAAD64646424B66E92241BAD6CDB64241C65659224ADDB246DB6B624),
    .INIT_1C(256'h1C8B1D1C93651B1B6C2424641B1BAD239292D21B1B24DB1C1CD3135C5D5D5C5C),
    .INIT_1D(256'hFDFEFEFEFEFEED6364F6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFFFFF658A),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDC41D36EF7FFFFFFFFFFB664EDEDF5F5F5),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_017408_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n28 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i17_008,inst_doa_i17_007,inst_doa_i17_006,inst_doa_i17_005,inst_doa_i17_004,inst_doa_i17_003,inst_doa_i17_002,inst_doa_i17_001,inst_doa_i17_000}));
  // address_offset=18432;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFE7FFFFFFFFFFE25F71B07FFFBFFFECFF86307FE0F3CFCFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFE25F61BFFFFFFFFBD9FF8E300610F78FCFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFC2BF61FFFFFFFFF7D9DF8E100000EF1FCFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFC2AE61FFFFEFFFEFB1FFBE1000005F3FCFFFFFFFF),
    .INIT_00(256'h6CF6FF646DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hA4A4641C641C1BDBD2DBDBDB1C241B1BD2DB6DB6AD2492DB246D6D24ADB5DADB),
    .INIT_02(256'h6C24D2DB6D6D641B6D246D6D24DBDBDBD364AD8A4B016D6D4A4B0A02931B64A4),
    .INIT_03(256'h1B5B5BA51B1BAD2364236DFFB69365AD1B2464246465651BAD232324B6B66CDB),
    .INIT_04(256'hD4D31DD4D365D264646464648964AD1B9191D21B1BDB1C1B8AD2D3D3D3131313),
    .INIT_05(256'hFEFEFEFEFEFEAC64F5F6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFFFFF248A),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDCDCAEF7FFFFFFFFFFFFFF64ADEDEDF5F5),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h24B6FF6D24FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hD31C2401014ADB23DBDBDBDB2424241BD26CB6B524DBDBDB6C6D1B24ADB5DBDA),
    .INIT_0A(256'h6DDBDA246D6C24246D246D6D24DBDBDB1C64AD934B01246D93035454535393D3),
    .INIT_0B(256'hACADAD5C5C1C646C1B641BF6FFB6646464646424656D24AE64DB24ADB66DDB24),
    .INIT_0C(256'hD4D31DD4DC24DB6C1C65642340AD6DD28991D21B1BDB1B2364A5ADADADADADAD),
    .INIT_0D(256'hF5F6FEFEFEFEFEF6F6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFFFFEFE1B8B),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF256EB7FFFFFFFFFFFFFFFF6D64F5F5F5F5),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h24B6FFFE24B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h9C939CDDE5E5DCDBDBDBDBDB242423DB24B6B624DBDADB24AD242424ADB6DBDB),
    .INIT_12(256'h24DBDB246D6CDB6C6C24AD6524DBDBDB66656DDB020A936D9B020B0B4B539493),
    .INIT_13(256'hF5F5ADEDA45B13646423636464A51C1B64641C2465656D6DDB246DB6B624DB64),
    .INIT_14(256'hD3D31DD31CDB64641C65641A89AD64D28991D21B1C1B63AC63A4A36363ACECF5),
    .INIT_15(256'hF6F6F6FEFEFEFEFEF6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFFFFFF589D3),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAEB7B7FFFFFFFFFFFFFFFFB624ACF5F5F5),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h246DFFFF6D6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h949CDDE5E6DCDBE3DBDBDADBDB24DB24B6B6241BDBDA2364AD242424ADB5DBDB),
    .INIT_1A(256'hDBDBDB6D64241B6D646D6D651CDB2425666D6CDB014B0125DC0A535353535394),
    .INIT_1B(256'hF5FEF5F5F5AD138A246C6C64EDEEEDAD246424656565AEDB2464ADB664DB2424),
    .INIT_1C(256'hD3D41DD31CDBADDB1C6564D1DAAD64918A92DA1B6463ACACABA3ABEBA2A3ECF4),
    .INIT_1D(256'hF5F5F5FEF6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFFEF65B41D3),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B7B7FFFFFFFFFFFFFFFFF7AE6CACF5F5),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_018432_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n28 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i18_008,inst_doa_i18_007,inst_doa_i18_006,inst_doa_i18_005,inst_doa_i18_004,inst_doa_i18_003,inst_doa_i18_002,inst_doa_i18_001,inst_doa_i18_000}));
  // address_offset=19456;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFBFFFFFFFC66EE3FFFFFEFFEF73FFFE000004BF3FCFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFE01FFFFFFFC66EC3FFFFFFFBDFF3BFFE08009C7B6FCFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFB407FFFFFFC64CC7FFFFFFFDBEE3BFFE00001CE4FFCFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFF003FFFFFFC6C8C7FFFFFEFF3EE3FFFF00000FB53FCFFFFFFFF),
    .INIT_00(256'h246DFFFFB624B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h9DDDDDE5E5DCDBDBDB23DADB23DB24B6B524246CDBDB6C1BAD6424246DB6DBDB),
    .INIT_02(256'hDB92246C6423246D6DAD6D242425252526AE24DB015301DCE44A5353949C949D),
    .INIT_03(256'hF5F5FEFDEDEDAD241BAD64D264EDEDED641B656565AE24DB246DB66DDB1B241B),
    .INIT_04(256'h8B1C1DD3D3246D8A24241B481BAD1B8989921B6464ACF4ECEBEBABABEBA2ABF4),
    .INIT_05(256'hF5F5F5F5FDFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFEFEFEF6A35B8A93),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6B7FFFFFFFFBFB7AE6E6D6565D3A4F5),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h246DF6FFFF246DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h9CDDE5E525DCDC241B1BDADADA64B66D23DB2424DB2424DBB62424246DB6DBDB),
    .INIT_0A(256'hDBD224246CDB6DB6256D65656D6D652525AE6D930A4B02931C4A0A0B4B539494),
    .INIT_0B(256'hF4F5FDFEF5ACADADAD1B1BB61B1BADA464D21B1CAE24DB246CB6B5231B242324),
    .INIT_0C(256'h8B1C1DD3D26D1C8A651C1B0064ADDB8989D2241B63ECF4F4F4F4ACABECEC63AB),
    .INIT_0D(256'hADF5F5F5F5F6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFEFEFEF563A4A400D4),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6B7FFFFB66D24DC8B8A8A01D48A415C),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h2424B6FFFF6D24FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hDDDDE5E5E59C9C252525DBDB6C6D64DBDB24DBDB231B2423B62424246DB6DBDB),
    .INIT_12(256'hD2DB246C24DB656D6D6D6E6E6E6E666E256EAEDC014B4B02DC930A4B4B539494),
    .INIT_13(256'hABF5FDFEFEFDF5F66D1BAD6D6D1BF6F6F6AD8A656DD324646DB624DB1B1B24DB),
    .INIT_14(256'h8B1D1D8AD26CD3D3251BDB0064ADD289891B641BACF4ECECECACACECACF5F463),
    .INIT_15(256'hD264F5F5F5F5F6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFEFEECA3A3F56341D4),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7B7B7B66E1CDB251CD41CD48B8B8A938A),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h2424B6FFFFB624B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h9D9DDDE5E59D01932525242464DB1B1BDB24921BDBDB241BB52424246DB6DBDB),
    .INIT_1A(256'hDADB242424246E6EAE6E6E6E6E6E6E6E6E6EAF6E014A4B4B52934A4B4B53949C),
    .INIT_1B(256'hABACF5FDFDF5FEF51BAD64D2646464F6F6AE656DDBDB246DB66D1BDB1B2424DB),
    .INIT_1C(256'hD31D1C8A2364D3D424DBD249ADAD9289881B2363ACACF4F4ECABACF4ECECF5F4),
    .INIT_1D(256'h82811BACF5F5F6F6FEFEFEFEFEFEFEFEFEFEFEFFFEFFFEFEACA3A3ECF51A4A8C),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7776E6EF7FFF7AE65D3D4D4D38B4A93D4),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_019456_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n28 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i19_008,inst_doa_i19_007,inst_doa_i19_006,inst_doa_i19_005,inst_doa_i19_004,inst_doa_i19_003,inst_doa_i19_002,inst_doa_i19_001,inst_doa_i19_000}));
  // address_offset=20480;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFC00FFFFFF84D8C7FFFFEDFF7CC7FFFF000007333FEFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFE103FFFFF84D9C7FFFFFF7EF9FFFFFF800007B33FEFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFF900FFFFF8CD9C7FFFFFFFFF1F1BFFF800007E77BEFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFF9003FFFF0DD9C7FFFFFFFFF39FEFFFC00003F77BEFFFFFFFF),
    .INIT_00(256'h24246DFFFFFF6D6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h949DDDE5DD9C0A93DC1C6D24DBDB2423DBDB1B64DBDB241BB52464246DB624DB),
    .INIT_02(256'hDA246D6EB7B7B6B6AEAFAEAE6E6E6E6E6E6E6EB7DC014B4B53534B4B4B4B9494),
    .INIT_03(256'hF4ACF5FDFEFEF6DAF5B5D21B1B641BF6FE6DAD1CDB246CB5AD24DBDB242C9AE3),
    .INIT_04(256'hD31DD48A641CD31C24DBD2D3AD6C8989481B2363ACEBECECECABACF4F4F4F4FD),
    .INIT_05(256'h8B8B42411CADF5F5F6FEFEFEFEFEFEFEFEFEFEFEFEFEEDA3A3A3E3F5F5928A8B),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6E6EB7FFFFFFFFFFFFAE24D3938B8AD3D3),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h24246DFFFFFFB624B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h9CDDE5DDDD4B4A94DC1CB6F76DDB2423DADB6C6DDBDB2423B52324246DB624DB),
    .INIT_0A(256'h6D76AEAEB6B7F7B7B6B6B6AEAE6EAEAEAF6E6EB76E014B4A4A939C9D9C949C9C),
    .INIT_0B(256'hFDF5ACF5FEFF64ADFEB41A1BD22423ADF66D23DB24656DB524DBDB1C651B236C),
    .INIT_0C(256'hD31DD4D3641BD31C24D3921CAD64888948232323ACABF4ECABECACECF4F4F4F5),
    .INIT_0D(256'h8B8B8B8A8A8A1BADF6F6FEFEFEFEFEFEFEFEFEFEF5A4A3E3E3E3ECF5AD498B8A),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B7FFFFFFFFFFFFFFFFB7B6DC4A4AD31C),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h24246CB6FFFFFF246DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hDDDDDD940B53DC9C9425AEFFF76D2492DB246D6D9A2364236DE324246CB6249A),
    .INIT_12(256'hDCDBDB1B1BD324F7B7B6B6B7B7B7B6AE6EAE6EB6B79C01530A0A4B949C9DDDDD),
    .INIT_13(256'hFEFEF5B5FEAD64FFFEAC1A1B1B1B6423B66C236D646DB66CDBDBDB6D6564AD64),
    .INIT_14(256'h131D93DB241BD31C24D2D21CAD63888A8823231BABABF4ABABF4ECACF4F4F4F4),
    .INIT_15(256'h938A8B8AD3CB418A1CADF6FEFEFEFEFEFEFEF6ECA3E3E3E3E3ECF5AD1C4A8A8A),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6FFFFFFFFFFFFFFFFFFFFFFB7258AD31C),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h2424246DFFFFFF6D64FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h534B4B4B9CE5E59C4BDCB7FFFFB62524DB246D6D9A2364246DDB246464B624DA),
    .INIT_1A(256'hA5F6FFFFFFF764DBFFB6B6B6B6B7B6B6B7B6AEB6B76E014B944A010A0A4B5353),
    .INIT_1B(256'hF5FEFEFEF523FEFFFEAC1B1A231B23246D6CB56C6CB6AD23DBDB6DAD24DBD21B),
    .INIT_1C(256'h1C1C931C1B1BD31C64D2DB1C6D63898A891B1B1BA3ABECABA3F4F4ECECF4F4F4),
    .INIT_1D(256'hD38A8B8AD3CB8B8B41411CADF6FEFEFEF6AD1AA4ECECECECACA4641C8A8A8A8A),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7FFFFFFFFFFFFFFFFFFFFFFB7B7D3D365),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_020480_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n36 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i20_008,inst_doa_i20_007,inst_doa_i20_006,inst_doa_i20_005,inst_doa_i20_004,inst_doa_i20_003,inst_doa_i20_002,inst_doa_i20_001,inst_doa_i20_000}));
  // address_offset=21504;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFF9000F1F0097BC7FFFFFFFFE7FFFFFFC00003FF7BEFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFF90000180097BC3FFFFFFFFCDFBFFFFE00003FF7BEFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFF7FF900000000B78C3FFFFFFFFFFFFFFFFE00083FFFBEFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFF07F980000000B78C3FFFFFFFFFFDFFFFFF78007FFFBE7FFFFFFF),
    .INIT_00(256'h24242424FFFFFFFF24B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h93949CDDDD9CE5940293B7FFFFB6FFFFB6246D6D92246424ADDB246424B664D2),
    .INIT_02(256'hDCEDF6FFFFFFFF1B6DFFB6B6B6B7B7B7B6B7B6B6F7B7940254944A094A4A9393),
    .INIT_03(256'hF4F5FEFE64ADFFFFFEF5631A631B64AD24FEAD24ADB524DBDA24AD651B6C6D64),
    .INIT_04(256'h1CDCD41CDA1B1C6565911B246D23488A891B1B1B63A3ECABA3ECF4F4ECECF4F4),
    .INIT_05(256'hD48B8B8A8BD38BCB8BCB8A8A1CAEAE6DDB0089EDEDAC6424DCDCDCDC8B8B8A8A),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6FFFFFFFFFFFFFFFFFFFFBFB7AF93D465),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h24242424B5FFFFFF6D6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h539394939CE5DD945393FFFFFFFFFFFFFFFFB66D92236C24ADDB246C24B66C9A),
    .INIT_0A(256'h12C112A5F7FFFFB61BFFFFF7F7F7B7B7B7B7B7B6F7FF66020B539C934A4A4B4B),
    .INIT_0B(256'hECB4FEF664FEFEFEFEFE641B23236DAD64F66D6DB66CDBDB2424D213ADFFFFAD),
    .INIT_0C(256'h1DD4DC24DA641C65AD891B1C6D23889289DB1B1B6362ECECA3ECF4F4F4ECACF4),
    .INIT_0D(256'hD4938B8A8AD3D38B8A8BD3D441418A00008A8A1C1CDB9393949C94534BD38A93),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6F7FFFFFFFFFFFFFFFFFFF76E8AD465),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h2364242464FFFFFFB624FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h534B94DD25DD94DD93DCFFFFFFFFFFFFFFFFFFFFB66D24246DDB236C24B66D9A),
    .INIT_12(256'hFFA54A019CFFFFFF1BB6FFFFFFFFFFB7B7B7B7B7B7FFB79C5394939C93535353),
    .INIT_13(256'hECF4FE64B5FFFEFEFEFEAC1B1B64646523AD6DADAD1B24B6AD1BADAD5C9CEEFF),
    .INIT_14(256'h1D8B2524DA641C65AD89DBDB6D23489289DA1B1B6362ECECA3ECF4F4F4F4ACAC),
    .INIT_15(256'hDCD38A938AD4D3D38A8A8BD3D38BD3D38A4A4A020A4B53535494DD9C4BD48AD3),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6D931C656EB6B6FFFFFFFFB7B76E41D466),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hDB64246C24FFFFFFFF6DB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h9CDDDDDDDD9CDDDD4B26FFFFFFFFFFFFFFFFFFFFFFFFB66D6DDB1B6C24B66DDB),
    .INIT_1A(256'hF6FFEE9301A4FFFF6C6DFFFFFFFFFFFFFFFFF7F7B7FFFF2D4AAEB66D25DC9393),
    .INIT_1B(256'hACF5AD64FEFFFEFEFDFEF51B2424236C63ADB6AE241BAEAE1BADFFFFEE53C19B),
    .INIT_1C(256'h1C8B6664D2AD1CAEAD89DBDB6D23489289D21B1B6362ABECA3ACF4F4F4F4ECAC),
    .INIT_1D(256'h1CD34A8B8B93D4D38A8A8AD3D38A8B8B8A4A0A0B5353949CDDDDDD948BD34ADC),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6938BDC8AD31C25B6FFFFB7B76542D466),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_021504_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n36 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i21_008,inst_doa_i21_007,inst_doa_i21_006,inst_doa_i21_005,inst_doa_i21_004,inst_doa_i21_003,inst_doa_i21_002,inst_doa_i21_001,inst_doa_i21_000}));
  // address_offset=22528;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFF3FF980000001B78C1FFFFFFFFFFF7FFFFF7F007FFFFE7FFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFF9C0000001778C1FFFFFFDFFFFB9FFFFBFC07FFFFE7FFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFDC0000041678C1FFFFFFDFFFFDDFFFF9FE07FFFF67FFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFEDC00000016F8C1FFFFFFDFFFFEFFFFFCFF0FFFFFEFFFFFFFF),
    .INIT_00(256'hDB6424641BB6FFFFFFB66DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hDCDCDDDDDDDD9C9D536EFFFFFFFFFFFFFFFFFFFFFFFFFFFFF61B136424AD6DDB),
    .INIT_02(256'hC1A4F7EE0A01A5FFB61BFFFFFFFFFFFFFFFFFFFFFFB7FFFF8A24FEFEF6B6AD24),
    .INIT_03(256'hACF563ACFEFEFEFEFEFEB5236C231B6463ACF6651C6DAD1CADAD64B5FEFFF613),
    .INIT_04(256'h1CD4AE64D2AD1CAEAD8993D36D2348D289D2DB1B6362ABF4ABABF4ECECF4F4F4),
    .INIT_05(256'h1CD48A8B8B8BD4D48B8A8A8BD38A8A8A8B4A4A4B5394949C9C9CDC8B93D44A1C),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7D3D32565AEB66D6D6EB6B7F76E42D4A6),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hDB246D242424FFFFFFFF6DB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hB66DDCDD9C949D9D94B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFF6125BAD1BADAEDB),
    .INIT_0A(256'hDC801BF6A5C1C1EEFF1CFEFFFFFFFFFFFFFFFFFFFFFFFFFF6D006DF6FEF6F6F6),
    .INIT_0B(256'hF5AD1BADF5FEFEFEFEFE6C64241BD2636C6CB6246D6D1BADAD6464636CB5FFFF),
    .INIT_0C(256'hD31DAE1CD2AD64B6AD498A936D6388D289D2DB1A63A3A3F4ABABF4ECACF4F4F5),
    .INIT_0D(256'h1D1C8B8B938A93D3D38A8A4A8AD3938A8B8B4A4A535393949CDDDC4ADCDC8A1D),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6656EB7FFFFFFFFFFB66E6EB7AED3D3AE),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hDB246D246C1BFFFFFFFFB66DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hF5FEB693539CDD9CDCBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9C01A5F6C1E5AD9B),
    .INIT_12(256'hF75B805BF7A5C152ED64B6FFFFFFFFFFFFFFFFFFFFFFFFFFBF939365F6F5F5F6),
    .INIT_13(256'hFE6463F5ACF5FEFEFEB564242463D16CAD64AD646D1B6DAD63ACF5F5F5B5ACB5),
    .INIT_14(256'h8B65AED2DAAD65F6AD8A4A8A646389D2D292DB1A63A3A3ECECABECECACACF4F5),
    .INIT_15(256'h1D1D8B8BD38A8AD3D38B8B8A8AD38B8BD4934A4B4B9494DDDD25D44ADC93931D),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B7F7FFFFFFFFFFFFFFB76E25AE2493AE),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h231B6D246D24B6FFFFFFFF6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hF5FEFF6E539DDD9425FFFFFFFFFFFFFFFFFFFFFFFFFFFFEE4A53EE640AEEF69B),
    .INIT_1A(256'h6DAE538064F7ED09A41BADFFFFFFFFFFFFFFFFFFFFFFFFFFFF6E018B1BACF5F5),
    .INIT_1B(256'hF61BADF5A3ABF5FEF624241B231BDAB5AD24AD6D1B65AD64ACF4F5FEFEFEFEB5),
    .INIT_1C(256'h8B6666411B6465F66D9392D364638992D292DB1A63A363ACF4ABECECECACACF5),
    .INIT_1D(256'h651DD38BD3D3938BD4938A8AD38B8BD4D34A4A4B539495DDDDDC938BDC53DC1C),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B7BFFFFFFFFFFFFFFFFFB7DCF7AE8A6E),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_022528_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n36 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i22_008,inst_doa_i22_007,inst_doa_i22_006,inst_doa_i22_005,inst_doa_i22_004,inst_doa_i22_003,inst_doa_i22_002,inst_doa_i22_001,inst_doa_i22_000}));
  // address_offset=23552;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFEDC002000067CC0FFFFFFFFFFFF7FFFFDFF8FFFF6EFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFEDE0060012C7CC0FFFFFFFFFFFFBFFFFFFF8FFFEFF7FFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFEFF0040002C7CC0FFFFEF7FFFFFDF7FFFFFCFFFEDFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFC6FBF890003C7860FFFF8FB83FFFFFFFFFFFEFFFF9FFFFFFFFF),
    .INIT_00(256'h1B236D646D6D6DFFFFFFFF6DB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hF5F5FEFF6DDCDD4B6EFFFFFFFFFFFFFFFFFFFFFFFFFFFF5CC1E5EEC1A4FFB6DB),
    .INIT_02(256'h6D6DAD0AC1A5FFF6A45B64F7FFFFFFFFFFFFFFFFFFFFFFFFFFB6D21B246423AC),
    .INIT_03(256'hAD1BFEF5AB63ACFEAD6D646DB52364B6B623B66524B664ACF4F5FEFEFEFDFEFE),
    .INIT_04(256'hD3AE6541DB6464AEAD1C93DC24649192D2D2DADA63A3A3ABF4ACECF4ECECACF5),
    .INIT_05(256'h6525D441D3D3D3D38BD393938B8B1CD442014B4B4B54949CDDDC8BD3DC4ADCD4),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6EB7FFFFFFFFFFFFFFFFFFB7DCB7F74A66),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hDB24646D246D24FFFFFFFFB66DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hABF5F6FFFFE493536EFFFFFFFFFFFFFFFFFFFFFFFFFFEDC113EE930AEEFEFE64),
    .INIT_0A(256'hFE6C6EAD0AC1A5FFFFA45B64ADFFFFFFFFFFFFFFFFF6F5ADADECF4F5F6FFF663),
    .INIT_0B(256'h6423FFFEF5ECEDADADADADF6F5ACB5F6B664F624F7ADACF4F5FEFEFEFEFEFEFE),
    .INIT_0C(256'h24AED441D3246464AE2501932364D289D2D2DAD263A3A3A3ECECECF4ECECACF5),
    .INIT_0D(256'h651C1D8A8A8B8BD3D3D4D48B8B1C1C4A4A4A4B4B4B4B539CE59C4A1DDC8B1DD3),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6DB6FFFFFFFFFFFFFFFFFFB793AEFFDB66),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h1B24246D246D6DB6FFFFFFFF6DB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hA4ACF5F5FEF69293B7FFFFFFFFFFFFFFFFFFFFFFFFF793C1E5A5C19CF6BEFFF6),
    .INIT_12(256'hFEFE6CAEEE53C19CFFB61BA4C19CF6FFFFFFFFF6B5F5F5F5F5F5F4F5F5FEFFFE),
    .INIT_13(256'h646DFFFEF6AC5BD212125B12D11A1B5B5B1A1B64F6ADF5F5F5FEFFFFFEFEFEFE),
    .INIT_14(256'h6D6E4A8BD31C2424B61C09931B64D289D2D2DAD25AA3A3A3ACECECF4ECECF4F5),
    .INIT_15(256'h651C6E65938B93D3D3D38B93D41C8A934B4A4A5393939CDDDD948BD44BD31DCB),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFB7B7B6B66EFFBF6DB7FFB7F7FFFFFFFFB7936DFF6525),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hAD24236D246D6D6DFFFFFFFFB66DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFEECECF5FEFFAEDCB6FFFFFFFFFFFFFFFFFFFFFFFFA501DCEECAC1EDF6BEFEFE),
    .INIT_1A(256'hBFFEF5ADB6EED341A46D6DEED40113ADFFFFFFFFF5EDF4F4ECF5F5F5F5F6FEFF),
    .INIT_1B(256'h24ADF6641A4080D1525A925A12D10A0A12C980D240D25B646363ADF6FFFFFEFE),
    .INIT_1C(256'hAE6501D3D31B6464B6DB4A49D2641B92D2D2DBD25AA3A3A3ABABACECF4ECF4F5),
    .INIT_1D(256'h65D46EFFAE251D1D66D48AD31CD38B1C4A4A530A4A539394938B8B4A01DC1414),
    .INIT_1E(256'hFFFFFFFFFFFFFFB7B66E6E6E6E256EFFB7B66D6E6E25DCDCDB256E9365FFF71D),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_023552_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n36 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i23_008,inst_doa_i23_007,inst_doa_i23_006,inst_doa_i23_005,inst_doa_i23_004,inst_doa_i23_003,inst_doa_i23_002,inst_doa_i23_001,inst_doa_i23_000}));
  // address_offset=24576;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFF0FBF88000587862FFFF3FE07FFFFFFFFFFFFFFFFBFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFB73F020005878E3FFFE7FE0FFFFFFF7FFFFFFFFBFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFF79E020003878E3FFFCFFFBFFFFFFFBFFBFFFFF77FFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFF7CC0600030F0D3FFF9FFFFFFFFFFBE7FFFFFFEEFFFFFFFFFF),
    .INIT_00(256'hFE6C1B6D6C6CB624FEFFFFFFFF6DBEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFEEDEDF5FEFEF5F5B6FEFFFFFFFFFFFFFFBFFFEE525BF6E4C15CB6B5FEFEFE),
    .INIT_02(256'hFEFEFEFEB5F5F6A55C5C64FFFF640941DBF6FFFFFFF6B6F6EDADADA4ADF5F6FE),
    .INIT_03(256'h5B5B5B12C9C912525A5A5A5A521209C98989C9D1D111115252525252ACF6FFFE),
    .INIT_04(256'hAED341D4D46565656E934A41D2241B91D2D21BD21AA3A3A2A3ABABECECF4F5F6),
    .INIT_05(256'h5DD465FFFFFFFFFFAE4AD3D41C82DCDC0A4B949C4B02024A4A8B93948B1CD31D),
    .INIT_06(256'hFFFFFFFFFFFF6EAEFFFFFFB7B66E76BFB7B76E76B66EAE1C0000DBD325FFFF25),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFEB5236C6D24B66DADFFFFFFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFEFEFEF5F5FEFEFEF6F6B6FFFFFFFFFFFFBFFFF653C1EEF60A53F66CB5FEF5FE),
    .INIT_0A(256'hFEFEFDFEFEF5F6F6F6645CADF6FFEE53C153E5F7FFFFFFFFF7F6F6B56464F6F5),
    .INIT_0B(256'h115B5BC9C9125A5A5A5A5A52521212C9898180C911125A9A9B9A9B5B125BF5FF),
    .INIT_0C(256'h6E418AD3D46E656D6D0101D3241B1BD2D2D21B1A5AABA3A2A2A3ABECECF5F6AC),
    .INIT_0D(256'hD4D41CFFFFFFFFFF8A4AD4D48B8B25DC024B4B949C945453938B934B931CD366),
    .INIT_0E(256'hFFFFFFFFB76DB7FFFFFFFFB76E6E6EB66E6EB7B6B6B7B7FFAE922425D3FFFFB6),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFEFE2423AD24B6B664FFFFFFFFFF6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFEFEFEFEFEFEFEFEFEFEADB6FFFFFFFFFFF7F69CC1E5F69BC9F6F66CB4F5FDFE),
    .INIT_12(256'hFFFEF5FEFEFFFEB5F6AD645C01E5F7FFA5C10194EEFFFFBFF7FFFFFFB6D264F5),
    .INIT_13(256'h125BC980529B9B9B5A5A5A5A5A52521212C91212125A529A9A9A9A9B5B5A5AED),
    .INIT_14(256'h2500D3D3DCAE646D250101DC6D1B1BDA92D1231A5AACABA2A2A3ABACF4F5AC5A),
    .INIT_15(256'h6541DB6EFFFFF7D30193D3D44ADC2593014B0A4A539494938A939493DCD41CAE),
    .INIT_16(256'hFFFFFFB7B6FFFFFFFFFFFFB66E6E252525B7B6FFB7B66EB7FFB6B66E8AF7FFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFEFE6C1BAD246DFF64FFFFFFFFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hF5FEFEFEFEFEFEFEFEFEFFB5B6FFFFFFFFF69CC05CF6E5C1EEF6ACF5ACB4FDFE),
    .INIT_1A(256'hADFEF5FEFEFEFFFEFE64ADF69BC15BEEF7EE9CC1CA5CAEF7F7B7F7FFFFAE12F4),
    .INIT_1B(256'h1180C95B9B9B9A5A5B9B9A9A5A5A5A5A52525B525A5B5A9A9A9B9A9A5A5B5A5A),
    .INIT_1C(256'hD342D38B1CAE646E93024BDCB7ADDB1BD2D1631A5AACABA3A2A3A3ACF5AC63A3),
    .INIT_1D(256'hFF65D3DC2465D3418BD3D38A932525934B4B4B4A02024A4B8B94DD94DCD365AE),
    .INIT_1E(256'hFFFFB7FFFFFFFFFFFFFF6E6E6E25252525FFB7FFFFB7FFB7B7B7F7B78AB6FFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_024576_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n44 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i24_008,inst_doa_i24_007,inst_doa_i24_006,inst_doa_i24_005,inst_doa_i24_004,inst_doa_i24_003,inst_doa_i24_002,inst_doa_i24_001,inst_doa_i24_000}));
  // address_offset=25600;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFF7F00600630F1F3FFF3FFFFFFFFFFEF1FFFFFFDDFFEFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFC0E00470F3F3FFE7FFFFFFFFFFF3CFFFFFF9BFFEFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFE1E00060F3F3FFFFFFFFFFFFFFFCFFFFFFFF7FFEFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFF3E00061E7FBFFFBFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hFEFE6CDB6D6D65FF6DB5FFFFFFFFFF6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hF5F5FEFEFEFEFEFEFEFEFEFFFEB6B6FFF7A4C052F6EDC1E4F6B5FDFDF4ACF5FE),
    .INIT_02(256'h5BACF6FEFEFEFEFEFE64B5F6F6ED0AC1DCEEF7ADC981C11365AD6EAEFFFFA4AC),
    .INIT_03(256'hC9C95BA39B9A9B9B9B9A9A5A5A9B5B5A5A9A5A525A5A9B5A9A5A9A9A5A9A9A9A),
    .INIT_04(256'h018B938B656D656D4A4BDC6DF7FF241BD2D1631A62ACECABA36363F5AC63A35B),
    .INIT_05(256'hFFFF651CDC4A018B8BD38B8ADC25254A0A535394949CDC938B1D2593DCD3AE6E),
    .INIT_06(256'hFFB7FFFFFFFFFFFFB66D6E6E2525B76E25FFFFFFFFFFB7FFFFB6FFFFD3AEFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFEFEADDA6D6D24FFB66DFFFFFFFFFF6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hF5F5F6FEFEFEFEFEFEFEFEFEFFFFFFF6AD81C1E5EE815BF6B5FEFEFDF5ECECF5),
    .INIT_0A(256'h9B9BACFEFEFEFEFEFE64FEFE75B6F6DCC1C1A4F6EE9CC1C91B6DAE6DADB5ACF5),
    .INIT_0B(256'h805BA35A5AA39B5A9B9A9A9A5A5A5A5A9A9A9A5A9A5A5A5A9A9A5A5A9A9A9A9A),
    .INIT_0C(256'h01938BD365656E254A5326B7B7FFB61BD2D2631A62ABACECA363ACACA3A35AC9),
    .INIT_0D(256'hAE6EAE6E6525D48A8B8A8ADC256E254B0A4B4B949DDDDD939425DCD4D31CAE1C),
    .INIT_0E(256'hB7FFFFF7FFFFFF6E6D6E6E256EB76E252DB7FFFFFFFFB6B7FF6EFFFF2465FFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFEFEF6DA24AD24B6FF6DFFFFFFFFFFB6B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFF6EECA13F6B5FEFEFEFEFEACACF5),
    .INIT_12(256'h9B9B9BACFEFFFEFEF564FFFFFFB6EDF6AE5C81C1A5EDE4ECF5FEFFFEFEFEFEFE),
    .INIT_13(256'h1B125A9AA35A529B9A9B9B9B5A525A9A5A5A5A5A9A9A5A5A5A5A5A9A5A9A9B9B),
    .INIT_14(256'h8B938BD36565AE254A94B7FFFFFFFF6DDAD2A35AA2ABACECECACAC63A35A0912),
    .INIT_15(256'h6E6EAEAE6E6525D48B8BD325656E254B0A4B4B539C9C948B94DC93DCD365AE8A),
    .INIT_16(256'hFFFFB7B7BFFFB66DB76F256E6E6EB66E2DB7FFFFFFFFF7B6B7B7FFFF6E1CAE6D),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6),
    .INIT_18(256'hFDFEFE1B23AD246DFF6DB6FFFFFFFFFF6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFEF6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFEDEEF6FEFFFFFEFEFEF5F5AC),
    .INIT_1A(256'h9B9B9B5BA4FEFFFFADADFFFFFFFEFEB56DEEE513C1A4ECECF4F5F5FEFEFEFEFD),
    .INIT_1B(256'h1BC95BA311119B9A9BA39B5A525A9A9A5A5A5A9A5A9A9A5A9B5A9A5A5A9A9BA3),
    .INIT_1C(256'h938B8A1C6666AFDC0125F7FFFFFFFFFF1BD2A35AA3ABECACECF5A49B5A0912A4),
    .INIT_1D(256'h6E6E6EAE6E252525D4421C256E6E25930A4B4B5354949393534A93D4D36E6541),
    .INIT_1E(256'hFFB7B6B6FFB76DB7B76E6E6EB76EB6B62DB6FFFFFFFFFF6E6EB6FFFF6E1C656E),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB76DB7),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_025600_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n44 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i25_008,inst_doa_i25_007,inst_doa_i25_006,inst_doa_i25_005,inst_doa_i25_004,inst_doa_i25_003,inst_doa_i25_002,inst_doa_i25_001,inst_doa_i25_000}));
  // address_offset=26624;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFF7FFF3E000C1E7FBFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFF7FFF3E000C1EFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFF7FFE7E00181CFFFFFF9FBFFFFFFEFFFF1FFFFFFFFFF7FFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFF7FFE7E00183DFFFFFB3F7FFFFFFEFFFFCFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hB5FEFE641BAD6D24FFB66DFFFFFFFFFF6DB6FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hF5F5F6F6FEFEFEFEFEFEFEFEFEFEFEFEF6AD5C9CDC9B9CEDEDF6F5FEFEFEFDB4),
    .INIT_02(256'hA39A9BA35B63FEFF64F6FFFFFEFEFEFEF5ADADADEDF5ECF4F5F5F5F5F5F5F5F5),
    .INIT_03(256'h12125BC9C99B9A9A9B9B5A125A9A9A9A9B5A5A5A9A9A9A9A9B9A9B9B5A9A9B9B),
    .INIT_04(256'h938B8B1D65AE6E01936EFFFFFFFFFFFF6CD1A362A3ABECACF5ED5B5A0912635A),
    .INIT_05(256'h6E6EAEAE65252525938B25256E6E25930B539354949393939353D4D31DAED38A),
    .INIT_06(256'hB7B66EB7FF6EB7B76EB7B66E6E6EFF766EB6FFFFFFFFFF6D936EB6B66E25256E),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6F7),
    .INIT_08(256'hB4FDFEADDA6D6D24FFFF6DFFFFFFFFFFB66DFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hECF5F5F6FEFEFEFEFEFDFEFEFEF6ED5B4A4A8B939293934A4A529BA4F5FEFEFD),
    .INIT_0A(256'hA39B9B9BA35A5BAD6DFEFFFEFEFEFEFEFEFEACF5F5ECF5EDA4A4A4A463A3ECEC),
    .INIT_0B(256'h5B1280C99B9B9B9B9B12115A9B9A9BA39B5A5A9B9B9A9A9A9A9B9B9A9B9A9B9B),
    .INIT_0C(256'hD38B8B6565AE250125B7FFFFFFFFFFFFAD1AABA3A3A3ECF4F5635209525B1212),
    .INIT_0D(256'hAE6EAE6E6565652541DC65256E6E65930A4B539494949394DC94D4D36E6641CB),
    .INIT_0E(256'h6E6EB7FFB6B6B76E6EB6B6B66EB7B76E6EB7FFFFFFFFFF6E0025B6B6B625656D),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6E),
    .INIT_10(256'hF5B5FEF6DA64AD24B6FF6DB6FFFFFFFFFF24FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hF5F5F5F5F6F6FEFEFEFEFEF6ED93014AD3D4D3939293D3D4D4D3D301A4FEFEFE),
    .INIT_12(256'h9B9B9A9A5BA45A88ADFFFEFEFEFEFEFEFEF5B4F5ECECA464D240CA1B1263F5F5),
    .INIT_13(256'h5AC9805BA39B9B9B12C95A9B9BA3A39B5252A39B5A9A9A9A5AA39B9B9B9A9B9B),
    .INIT_14(256'hCB8BD36565B7DC93B6FFFFFFFFFFFFFFF61AABA3A3A3ACF5AC1212525A12125B),
    .INIT_15(256'h6EAEAE6E6E6D6EDC4A2525656E6E65930A4B0B4B939393DCDD94D31CAEDC8AD3),
    .INIT_16(256'h6EB7B7B7B66E6E6E6D6EFFFFB6FFB66DB7B7FFFFFFB7FF6E926EB7B6B66D6565),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB724),
    .INIT_18(256'hFEB5F6FE2324AD6C6DFFB66DFFFFFFFFFF6DB6FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hF5F5F5F5F5F5FEF6FEFEED9C424293D48B424A935B93534A01014A015BFEFEFE),
    .INIT_1A(256'h9B9B5A9B5A9B9BC912ADFFFFFEFEFEFEFEFEECA3ACACAC6C641B814064F6F5F5),
    .INIT_1B(256'hC94012A39B9B9B12C95BA39B9B9B5B5252A3A35A9B5A5A9B5A9B9B9B9B9B5A9B),
    .INIT_1C(256'hD38A1C6565AE4A25B7FFFFFFFFFFFFFFF663ABA3A3ABADF55B11121212C95B5A),
    .INIT_1D(256'h6EB7AEAE6EAE6E8ADC25656E6EB66ED34B535494DC9394DDDCD493656E8A8B8B),
    .INIT_1E(256'h6EB7B7766E6EB66EB6FFFF6E6EB76E6DB7B7F7F7BFB6B7B6D3AEB6B6B6AE6E6D),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2D6E),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_026624_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n44 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i26_008,inst_doa_i26_007,inst_doa_i26_006,inst_doa_i26_005,inst_doa_i26_004,inst_doa_i26_003,inst_doa_i26_002,inst_doa_i26_001,inst_doa_i26_000}));
  // address_offset=27648;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFF7FFEFE00183DFFFFE67EFFFFFFFFBFFFFFFFFFFFE7FBFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFDFE00303FFFFFCC7DFBFFFFFFDFFFFFFFFFFFFFFFFFDFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFBFF9FE00303FFFFE08FBF7FFFFFFEFFFFE7FFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFBFF3FE00603FFFFE18F3CEEFFFFFF7FFFF03FFFFF7FFFFFFFF),
    .INIT_00(256'hFEFEB5FE6CDBAD6D6CFFFF6DFFFFFFFFFFB624FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hF5F5F5F5F5F5F5F6F5A452418BD34A015BEDF7F7FFFFF7F6F6A55C8189FEFFFE),
    .INIT_02(256'h9B9B5A5A9B5A5A5212C9ACFFFFFEFEFEFFFEFDECACACACACAC641B64F6F5F4F5),
    .INIT_03(256'h80095B5A5A9B12805BA39A9A9B5B1212A3A3529B5A5A5A5A5A5BA35B5A9B5A5A),
    .INIT_04(256'hD38A1C65AE65D36EFFFFFFFFFFFFFFFFFE64ACABA3ACF5AC121112D2C9525BC9),
    .INIT_05(256'h6EB7AEB6AEB61C4A25656E6E6EB76EDC025354949494939494D3D3AE1C8A8BD3),
    .INIT_06(256'h2576B66D76B7B7B6B7FFB7B66DFFB76E6EB7B7B7B776B7B7D365F7B6B6B6AE6D),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB66DB6),
    .INIT_08(256'hFEFEFEFEF51B6DAD24FFFF6DB6FFFFFFFFB6DBFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h5B64A4ACEDF5F5EC524A92938A0153EDFFFFF7F6EDEDEEF6F7F7F6EE64F6FFFE),
    .INIT_0A(256'h9B9B5B529B5A11A35212C9ACFFFFFEFEFEFEFEFEFDF5ACABABA3A4EDF5ECEC63),
    .INIT_0B(256'h805B9B125B12405BA45A9AA352C912A3A3125B9B125B5A5A5A5AA35A5AA39B52),
    .INIT_0C(256'h8B8B1D65AE1C25B7FFFFFFFFFFFFFFFFFF6CACABABACF55B1111D189125BC980),
    .INIT_0D(256'h65AEB7B6F76E011C6E6D6EAEB6B76EDC010B4B4A93934B94D48B656E8B8B8BD3),
    .INIT_0E(256'h6E252D6EFFB7FFB7B6B76EB7B7FFB76E6DB6B7B7B66EB7B7131BF6B6B7B7B66E),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7B7B7B6FF),
    .INIT_10(256'hFEFEFEF5FE6464B564B6FFB66DFFFFFFFFFF246DFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h40131B1364A49C529393930152EDF7F7EEA4534A4A4A4A52539CA4E5ADF6FFFE),
    .INIT_12(256'h5AA35A12525A529B5B521280ADFFFFFEFEFEFEFEFEFEFEF5F5ECACECECEC6340),
    .INIT_13(256'h12A4125B12401AA45A5BA312C85AA3A3115AA312129B115A525AA35B529BA35A),
    .INIT_14(256'h8AD31D65AE256EFFFFFFFFFFFFFFFFFFFFACACABACF5A4D1D1D189C95BD2C180),
    .INIT_15(256'h6D6EF7F7AE8BD3AE6E6EB7B6B6B7AEDC014B4B4B939394DC93D36E1D8A8BD3D4),
    .INIT_16(256'hBF25B7FFB7FFFFB6FFB76E6EFFFFB66E6EB7B7B7B7B6B7F75CC1AEB7B7F7B7AE),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6FFB7B7FF),
    .INIT_18(256'hFEFEFEFEF56C23B565ADFFFF6DFFFFFFFFFF6D24FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hD3418BD38ACA5393D38B4AE5F7F7AD1B018ACBCBCBCBCBCBCB8B4A4ACA64FEFE),
    .INIT_1A(256'h11A39A52115B5B5A5B12520A80ADFEFEFEFEFEFEFEFEFEFEFFF6ECECECA45C1C),
    .INIT_1B(256'h635B121240D2A45A5A5BC9C95B9B9BC9529B5AC95B5A095B5252A39B529BA35A),
    .INIT_1C(256'h8AD41DA66E65B7FFFFFFFFFFFFFFFFFFFEACECABECEC1AC9D189801212C980C9),
    .INIT_1D(256'hAE246DAED341AEAF6EB7B7B6B7F7AEDC02535393D393DC948B1C6ED38B8BD3D4),
    .INIT_1E(256'hFFB6FFFFB7B76EFFFFB725B7FFFFB66E76B7B7B6F7FFFFF7A58165BFBFF7F7B7),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6FFFFB7B7BFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_027648_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n44 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i27_008,inst_doa_i27_007,inst_doa_i27_006,inst_doa_i27_005,inst_doa_i27_004,inst_doa_i27_003,inst_doa_i27_002,inst_doa_i27_001,inst_doa_i27_000}));
  // address_offset=28672;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFDFE7FE00603FFFFC11E79DDFFFFFF3FFFFCFFFFFFFFFFFEFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFDFFFFF00C23FFFF801EF39DF7FFFF9FFFFEFF7FFFFFFFFEFFF),
    .INITP_02(256'hFFFFFFFFFFFFC0FFFFFF00C27FFFF803CC73BB7FF7F9FFFFCFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFC16FFFFF00867FFFF00380F7337FF7F8FFFFE7FFFFFFFFFFFFFF),
    .INIT_00(256'hFEFEFEFEFEB423AD6D6DFFFF6DB6FFFFFFFFB6DBFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h641CD2814A93D3934A5CF6FFEE9341824A4A525B5B5C5B531352528A4201EDFE),
    .INIT_02(256'h119B9B09115A9B525B5A1212C980EDFFFEFEFEFEFEFEFEFEFEF5ECECABACACA3),
    .INIT_03(256'h9B125BC989A35A5A5B81C95B9B5BC9125B5BC9125B51095B1212A39B125BA3A2),
    .INIT_04(256'h8AD41D6E656EF7F7F7FFFFFFFFFFFFFFFEACECACF5A480CA89808912C989801A),
    .INIT_05(256'hF7AE1C418AAEF76EB6FFFFB7B7B7B6DC025353949394DC9393651D4A9393DCD3),
    .INIT_06(256'hFFBFFFFFB6B6FFFFFFB6B6FFFFBF6E6EB7B7B7B6B777776E6D13CAEEFFBFFFF7),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7FFB7FFFFB7FF),
    .INIT_08(256'hFEFEFEFEFEFE236DAD64FFFFB66EFFFFFFFFB6DBB6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h646464CA53934A53EEF7F69CC14A4A0153A5F6FFFFFFFFF7F6F6EDE5DD535CFE),
    .INIT_0A(256'h119B9B0909525B5B525B12121289C9F6FFFEF5B5F5FEFEFEFEF5F5ACABACA3A3),
    .INIT_0B(256'h5A1212405B5A121280C9535B5BC9C95B5B11C95B5A11115BC9129B9B115A9BA3),
    .INIT_0C(256'h8BDC65AE65B6F7F7FFFFFFFFFFFFFFFFFEACECF5F5D2C9C98180C9C9C989C95B),
    .INIT_0D(256'hFFFFF76EB6FFB7AEB7FFFFF7FFFFB7240A53939C93DCD48B1C65D38B8BD31C93),
    .INIT_0E(256'hFFFFFFB6B6FFFFFFB7B7FFFFFFB66D252D6EAE651C1C2565ADA5C19CFFFFBFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7FFFFFFB7FFFF),
    .INIT_10(256'hFEFEFEFEFEFEB524B624B6FFFF6DFFFFFFFFFF236DFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hF56CD281020A64F7FFE50A4A4B0253ADF7FFFFFFFFFFFFFFFFFFFFFFFFF7ADB6),
    .INIT_12(256'h115A9B09C9525A5B525A521212C9401AF6B5ADFEFEFEFEFEF6B5ACABACACACF5),
    .INIT_13(256'h121280D21211C980C952525AD1885A5A1280125B12C9125AC9129B5B111A5B9B),
    .INIT_14(256'h931C65666EB7B7FFFFFFFFFFFFFFFFFFF6B5F5F56440D1C98980C9C9C9C9125B),
    .INIT_15(256'hFFFFFFFFFFFFB6B7FFFFFFFFFFFFB7250B93939393DC948B651D42938BD41C8B),
    .INIT_16(256'hFFB7B7B6FFFFFFB7FF6DFFFFFFFFBFB66E1C8A8AD38A41811BE59301F6FFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFEFEFEFEFDFEFEB5B56DB6FFFFADB6FFFFFFFF246DFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFEF51A404113F6F75C014A420BA5F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBE),
    .INIT_1A(256'h12129B11C912525B5252521112C9C98063FEFEFEFEFEFEFEFEF5B4F5F5F5FEFE),
    .INIT_1B(256'h12C988D1C9C988C91212121180125B1289C95A52D28912128012A45A11125A9B),
    .INIT_1C(256'hD31CA665AEB7B7FFFFFFFFFFFFFFFFFFF5B5F5F588C9D1C98081C9C9C9C95252),
    .INIT_1D(256'hFFFFFFFFFFFFB7BFFFFFFFFFFFFFB7250A93949393DC8BD465D38AD3931C1C8A),
    .INIT_1E(256'hB7FFB7B7FFFFB7B6B66DFFFFFFFFFFFFFF1C42CBD48AD35CC9E4E5C19CFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6FFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_028672_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n52 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i28_008,inst_doa_i28_007,inst_doa_i28_006,inst_doa_i28_005,inst_doa_i28_004,inst_doa_i28_003,inst_doa_i28_002,inst_doa_i28_001,inst_doa_i28_000}));
  // address_offset=29696;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFDBF7FFFF01847FFFF003018E727FF7FA7FFFEEFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFD3BFFFFF01047FFFE403000C627FE7FB7FFFF87FFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFF3DBFFFF030C7FFFE4060008C06BE7F9BFFFF8FFFFFFFFFFF7FF),
    .INITP_03(256'hFFFFFFFFFFFFF7FDFFFF020CFFFFEC2008628863E7F5BFFFF9FFFFFFFFFFF7FF),
    .INIT_00(256'hFEFEFEFEF5F5FEFEB56C6DFFFFF66DFFFFFFFF6D24FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFEFD63891C251C814A93025CAEF7FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'h12125B11C812525B5A115A0912C91BD2C9F6FFFEF5FEFEFEFEFEFEFEFEFEFEFE),
    .INIT_03(256'hD28989C9C981801212D2D288095212C98812521289C912D28012A4120912529B),
    .INIT_04(256'hD31C6665B7B7B7FFFFFFFFFFFFFFFFFFB5F5F61B40C9D1C98989C9C9C9C95A12),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7654B4BD49394948A651D41D38BD31DDC8A),
    .INIT_06(256'hFFB6B6FFFFFFB7B76DFFFFFFFFFFF725F7AE8A1D1C001CF65253ED5CC1EDFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7FFFF),
    .INIT_08(256'hFEFEFEFEFEF5F5FEFE6C6CFFFFFF6DFFFFFFFF6D24FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFDAB1A64DB40C1C153EEF7B6B6B7FFFFFFFFFFFFFFFFFFF7F7FFFFFFFFFFFF),
    .INIT_0A(256'h12125BC9C812525A5A11521212C95B64801BFEFEF5FEFEFEFEFEFEFEFEFEFEFE),
    .INIT_0B(256'h898189898180C9C9C9C989C91212C9C9C91212C989D112CA8912A3111112525A),
    .INIT_0C(256'hD365656EB7B7B7FFFFFFFFFFFFFFFFFFF5FEAC80C912D1898989C9C9C9D21211),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6E4A4AD38BD48BD365D342D38AD41DD48A),
    .INIT_0E(256'hB6B6FFFFFFFFB7B6B6FFFFB7FFFFB66DFFB7DC65D3001BF6EDC1A5ED5293F7FF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7B6),
    .INIT_10(256'hFFFEFEFEFEFEB4F5FEF524FEFFFFB5B6FFFFFFB5DBB6FFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFEAB621B40898113ADFFFFFFB6B6F7FFFFFFFFFFFFFFFFF7F7F7FFFFFFFFFF),
    .INIT_12(256'h12125AC9C912125A5A12125209CAD2B612C9B5FEF5FEFEFEFEFEFEFEFEFEFEFE),
    .INIT_13(256'h8989898989C9C9C9C9C9D2D212C1C9C91212C980D2D2C9C989125BC911C9525A),
    .INIT_14(256'hD46565AEB7B7FFFFFFFFFFFFFFFFFFFFF6F51AC9C912C9C980C9CAD2C91212C9),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6E4A4B938B944A1D1D418B938B1C1DD38B),
    .INIT_16(256'hFFFFFFFFFFFFFFAEFFFFFFF7FFFFF76EFFB724658A8A23ACF65CCAEDDCC15CFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B7),
    .INIT_18(256'hFFF6FEFEFEFEF5ACF5FEADB5FFFFB66DFFFFFFB6DBB6FFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFEF4621A40811C6E76B6FFFFFFB6B6FFFFFFFFFFFFFFFFFFF7F7FFFFFFFFFF),
    .INIT_1A(256'h111112C9C912125A5B111252C91240B6A48063F6F5F5FDFDFEFEFEFEFEFEFEFE),
    .INIT_1B(256'h898980C912C9C9D2C91A12D281C912D212D180C912C9D2D2891212C9D1C9125A),
    .INIT_1C(256'h1C6565B6B7B7FFFFFFFFFFFFFFFFFFFFF6631AC91212C9D1C9C912C9C9C9C9C9),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAE4A9393938B9325D341D48BD31C5D8B93),
    .INIT_1E(256'hFFFFFFFFFFFFB7FFFFFFFFB7B7FFB71C6EB6241C0112A3ABF6EE01DBEE1381E5),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_029696_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n52 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i29_008,inst_doa_i29_007,inst_doa_i29_006,inst_doa_i29_005,inst_doa_i29_004,inst_doa_i29_003,inst_doa_i29_002,inst_doa_i29_001,inst_doa_i29_000}));
  // address_offset=30720;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFE7FDFFFF060CFFFFF8E412C61B4367F1BFFFFBFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFE7F6FFFF041CFFFFDB45B7CC134347F1FFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFF4FF67FFF8418FFFFB3516F98364307D1DFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFE4FFB3FFF8C19FFFF73D3433966D207D1DFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h646CFEFEFEFEFEACABFDFE6DFFFFFF6DFFFFFFB61BB6FFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFEFEF5635B891C666E6EB6B6FFFFFFFFFFFFFFFFFFFFFEF6B5ADACACA463ACAD),
    .INIT_02(256'hC91212C9C912125A5B121152C9D240ADED801BF5F5F5F5F5FDFEFEFEFEFEFEFE),
    .INIT_03(256'hD280C912C9C912C95B5BC980895B12CAD280801212401A12C952C988C9C91252),
    .INIT_04(256'h1D6566B6B6F7FFFFFFFFFFFFFFFFFFFFA31A12095BC9C9CA120912C9C912D1C9),
    .INIT_05(256'hF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFB6D38B938B4A1C1D418BD48BD4251D8AD3),
    .INIT_06(256'hFFFFFFFFFFB76EB6FFFFFFB7B7B61CB6BF651C94015BA3A3ADF69C01E5A58149),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hF66CFDFEFEFFFEF563F4FE6CFFFFFF6DB6FFFFB624B6FFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFEFEF563631B65666EAEB6B7FFFFFFFFFFFFFFF6AD646463ACF5ECA35AABFDFE),
    .INIT_0A(256'hC912C988C912095A5A120952C9D14064ED1212ADF5F5F5F5F5F5F5FEFEFEFEFE),
    .INIT_0B(256'h12405B12C95B125BAC128080A46389CA8980C95BC9895B11C85BC9C988C91212),
    .INIT_0C(256'h1D656EB7B7F7FFFFFFFFFFFFFFFFFFA4125AC95B12C91209C912C9C9C912C912),
    .INIT_0D(256'h5CF7FFFFFFFFFFFFFFFFFFFFFFFFFFB6DC8B8B4A8B1DD401D3D38B1C651C8AD4),
    .INIT_0E(256'hFFFFFFFFB6FFB66DFFFFFFB7B6B6B6F76E1C1D8A8A63A3ABACF5ED0AC1E65CC0),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFF5ACFDFEFEFEFEACACF56CFFFFFFB66DFFFFAD24B6FFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFEFEFDA3636425256E6EB6B7B7FFFFFFFFF66C63A3A3ACF5FEFDECA3F4FEFEFF),
    .INIT_12(256'hC9CAC989C912115B1A12C912C9C94064EDA3C9ACF5F5F4F4F5F5F5F5FDFDFEFE),
    .INIT_13(256'h88126480636363ED634088ECECC9C9C9C9C9A35B0063A4C8C912C9C9C9C91212),
    .INIT_14(256'h6565AEB7B7FFFFFFFFFFFFFFFFFFA4125AC95A5BC9C9520AC912C912C9C9C95B),
    .INIT_15(256'hC1A5FFFFFFFFFFFFFFFFFFFFFFFFFFFF1C8A8B4AD41D8A8AD38B8B1D65DC8BD4),
    .INIT_16(256'hFFFFFFFFB6246EFFFFFFFFB7B66EB765D31DD4411BABABA3ACACFEA58152EDD3),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFEF5ACF4FEFEFEFEFDACAC64B6FFFFFF65FFFF6D24FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFEFEF5626364252E6E6EB7B7B7FFFFFFAD6363EBEBF4F5FEFEF56BB4FEFEFFFF),
    .INIT_1A(256'hC9C980C9C912125B1212C912C9C94064A3ACD1A4F5F4F4F4F4F5F5F5F5FDFEFE),
    .INIT_1B(256'h891BD200D1D2ADAD40C9ACF512408012C95BAC89D1ADA380121BC912C9C912C9),
    .INIT_1C(256'h6525B6B7B7FFFFFFFFFFFFFFFF641212C952A312C9C90A520A12C912C9C91264),
    .INIT_1D(256'hC1C1ADFFFFFFFFFFFFFFFFFFFFFFFFFF1D8A8B4A1C1C418BD38AD36566D39314),
    .INIT_1E(256'hFFFFFFB6F7F7B7FFFFFFFFB76E256EDBD4668B81A3ABABA3ABACB5F612805C6E),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_030720_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n52 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i30_008,inst_doa_i30_007,inst_doa_i30_006,inst_doa_i30_005,inst_doa_i30_004,inst_doa_i30_003,inst_doa_i30_002,inst_doa_i30_001,inst_doa_i30_000}));
  // address_offset=31744;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFCFF9BFFF0819FFFFE9D30073EED00B95FFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFF9FFCDFFF1839FFFFF07201E7DC300B57FFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFDFFF9FFE6FFF1039FFEFF01603CFD80007E7FFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFF90FFBFFE77FF10397FDFF0E403FFF80406EF7FFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hFEACECF4F5FEFEFEFEB56464B6FFFFFF6DFFFF6D64FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFDFEEC62A36324666E6E76B7F7FFF66362A3ECECF4FDFEFEFD6CB5FEFEFEFEFE),
    .INIT_02(256'hC98989C912C9525B12D2C9128012D2645AEC1A63F5F4F4F4F4F4F4F4F5F5F5FE),
    .INIT_03(256'h008940400000DAD2D2ADF6A440405B1B5BF56300ADF51280121AD15B80C9D2C9),
    .INIT_04(256'h2525B7B7F7F7FFFFFFFFFFFFA412121212A45BC912C9C0090A12C91289C9645B),
    .INIT_05(256'hA48112F6FFFFFFFFFFFFFFFFFFFFFFFFDC8A4A93258B8A8BD38AD4666693D31D),
    .INIT_06(256'hFFFFF76DF7AEFFFFFFFFBFB76D256E256E2541D2ABABABA362ACACADA58181A5),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hF5ACACF4F4F5FEFEFEFEAC6CADFFFFFFB6B6FF6D6DFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFDF5ABABAB6364656E6EB6B6B6AC6262A2EBACF5FEFEFEFEACB5FEFEFEFEFEFE),
    .INIT_0A(256'h8980C9C912C95B12D212D212805B1B645AAC6363F5ECF4ECF4F4F4F4F4F5F5F5),
    .INIT_0B(256'h004880884049891BEDF6AD4089A4A463F5F5D21BF61A40C989401B1B40CAC989),
    .INIT_0C(256'h2425F7B7F7F7FFFFFFFFFF6411121212A3A31112D1C980C9C90A0A1288D164D2),
    .INIT_0D(256'h655CC153F7FFFFFFFFFFFFFFFFFFFFFFD38A421C1C8A8AD3938A1CAE658AD31D),
    .INIT_0E(256'hFFFF1C65F7AEFFFFFFFFB7B625256E6EAED34164ABABABA362ABF4A4AD5C80C9),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hB4F5ECF4F4F5FDFEFEFEF56C6DFFFFFFB66DB66D6DFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hF5F563ECABA364646DAEAD6D635AA3ACF4F5FEFEFEFEFEF5B4FEFEFEFEFEFEFD),
    .INIT_12(256'h818189C9C9125B12121B12C989AC646308A36463F5ECECABF4ACACF4F4F4F5F5),
    .INIT_13(256'h49488080490024F6F6F5D1D2EDF5A4F5F6ACDAB5240089894000D2D180C9C981),
    .INIT_14(256'h1C6DB7B7B7B7FFFFFFFFA4C95B5B529BA3520A12C980818080C9C10A801A1B89),
    .INIT_15(256'hD2A55BC15CF7FFFFFFFFFFFFFFFFFFB68B8A8A1CD38B8BD38B931DAE658AD365),
    .INIT_16(256'hFFB6011DAEF7B7B6FFFFB725B66E25AE6641D2ACABABABA363ECF4F4646D1380),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hF5FEFDACF5F5FDFEFEFFFE6C6CFFFFFFFF246D6DADFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hF5AC63F4E3A3636C6D6D65A4ECF4F5FEFEFEFFFEFEFDF4ACFEFEF5FEFEFEFEF5),
    .INIT_1A(256'h8189C9C9C95B5BD212A412401BAD645BC05B646CF5ECABF4F4ACACF4F4F4F4F4),
    .INIT_1B(256'h0040894089006DFEF66363F5F6EDF5FDF6ACACFEADD2408980890040D2128081),
    .INIT_1C(256'hDB6DB7B7B7F7FFFFFFADC05BAC1A5BDB5A111212898980C9645B0AC18023DA00),
    .INIT_1D(256'h4013AD9CC19CFFFFFFFFFFFFFFFFFF6E8A42D41C8B8BD3D38AD465AE1C8BD465),
    .INIT_1E(256'hFFD38B1CD3414A9324B6B725B6B665AF154163ACABABA3A3A3EDF5F4AC6365D3),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_031744_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n52 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i31_008,inst_doa_i31_007,inst_doa_i31_006,inst_doa_i31_005,inst_doa_i31_004,inst_doa_i31_003,inst_doa_i31_002,inst_doa_i31_001,inst_doa_i31_000}));
  // address_offset=32768;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFB01F3FFF3FFF207BFFFFE1E4C3FFF8080ECF7FFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFF22477FFF9DFF2073FFB7C1FF83FFFE0006DF7FFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFF42EE7FFFE07F4073FFFF81FF8BFFFE040DDEFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFEC4DEFFFFE37E4073FFFF01FEDFFFFE0C1BBFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hFEFFFEF5F5F5FDFEFEFEFEF564FEFFFFFF6D246DB6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hF4ABA3F4AB63636362A3ECF5F5F5F5F5F5F5F5F5F4ACB4FDFDB5FEFEFEFEF5FE),
    .INIT_02(256'h8989C9C9125B9C406CB5C980ADB52311C05BACACF5ACACF4ECABECECECF4ECF4),
    .INIT_03(256'h641A4081C940B5FEF5F5F6F6F5F6F5F6F5F5FDFEB5004088808088881AD14081),
    .INIT_04(256'h1CAEF7F7F7B7FFFFFE1A23F65B51A363121212C989C9401BF563ACD1C91BD2DB),
    .INIT_05(256'hCA401BF6E5019CF7FFFFBFFFFFFFFF6D418A1CD38B8BD4D38A1C65AF1C8A1C65),
    .INIT_06(256'h66411D1DD48BD38B0141D466AF656E6E8AD3ACACECABA262A3F5F5F5FDAC6464),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFEFEFEB5FEFDFDFEFEFEFE6CB6FFFFFFB66D6DB6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hF4A3ABF4AB63A3636263A3A3ABABACACACECACACACF4F5F4ACF5FEFEFEFEFEFE),
    .INIT_0A(256'h8981C9D289AD5B81B6AD4012F6AD1B09C063ACACF4A3ECF4ABABECF4F4F4F4F4),
    .INIT_0B(256'hFEDA40D28940F5FEF6F6FEF6FEF5F5FEF6F6F6FE6D64644080404189D188C989),
    .INIT_0C(256'h24B6B7B6B7BFBFFFADD2F6ADC99BA35A5252C98989C90064F563EDA312AD6CB6),
    .INIT_0D(256'h1CD38A64ED5BC95BF7FFFFFFFFFFFF2501D41C8BD38BD48B8B1DAEAFD38B1D65),
    .INIT_0E(256'h8AD41DD4D38B1CD3DC1C8BD3DC25AF1C4164ACECEBA3A362ACF5F5F5FDF66464),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7),
    .INIT_10(256'hFEFEFEFEF5F5FEFEFEFEFEFFB5B5FFFFFFB66D6DFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hAC63ABF4ABA3A3A3A362ABABABABABABABACABECF4F4AB63F5FEFEFEFEFEFEFE),
    .INIT_12(256'h89C9C940ADAD4064F61B40A4EDAD5B8010ABF5F4ABACF4ACAAABECF4ACF4F4F4),
    .INIT_13(256'hF5DA00D26489F6FEFEFEFEFEFEFEFEFEFEF6FEFEADF7AD40898941928912D2C9),
    .INIT_14(256'h25B6B7B6B7FFFFFF1BADF6125AA39A5A52C9C98989894064F5ACECEC1AF5B56D),
    .INIT_15(256'h242423DBDBD2D2D2DBB6FFFFFFFFFF24011CD48BD38BD48AD365AEAE93D3651D),
    .INIT_16(256'h931DD4D38BD41C8B1C1D1CDC24AEAE8BD2ACECECABA3A262F4FEF5B5AC6C2424),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1C),
    .INIT_18(256'hFEFEFEFEFEB4F5FEFEFEFEFEFEB6FFFFFF6C6DB5FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hAC63ECECABA2A2A3A3A2A3ABABABACF4F4F4ECECAB6363F5FEFEFEFEFEFEFEFE),
    .INIT_1A(256'hC98088ADFF911BA4ADD21AECA4A35A11A2EBACACA3ACF5ACABACECF5F4F4F4F4),
    .INIT_1B(256'h1A638811AC64FEFEFEFEFEFEFEFEFEFEFEFEFEFE64641B40C98949D31B12C9D2),
    .INIT_1C(256'h25AEF7F7F7EEEDAD1BF66412A39B5A52C9C9898989CA401BF5ECA3ECA3F5F5DA),
    .INIT_1D(256'h232324DBDBDB1B23DB1B6DAEB6FFFFDB421D8BD3D3D3D441D465B6AE8BD4651D),
    .INIT_1E(256'h1C1CD48B8B1CD4D31C1DD465AEF71C4263ACECECABA363ABF5B56C232323231B),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAE41),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_032768_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n60 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i32_008,inst_doa_i32_007,inst_doa_i32_006,inst_doa_i32_005,inst_doa_i32_004,inst_doa_i32_003,inst_doa_i32_002,inst_doa_i32_001,inst_doa_i32_000}));
  // address_offset=33792;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFC84BCFFEFDBFE40F7FFFE01FF73FFFE967FFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFD0CBDFFFFFFFF80F78FFC00FF43FFF7BCFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFA097BFFFFF38F84F79FF8007F7FFFFBF9FFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFF8197BFFFE207EC0F7FFF3003FFFFFFE7E7FFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hFEFEFEFEFEFDACF5FDFEFEFEFFFEFFFFB66D6DB6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hABA3ECECABA2A2A2A3A262A2A3ABACECECECABA363ACFDFEFEFEFEFEFEFEFEFE),
    .INIT_02(256'h401BB5FF1B1BAC636412A49A599A62A2A3A3ACA3ADF6F6F6EDEDEDF4F4F4F4F4),
    .INIT_03(256'h80ECEB5A88DABEFEFEFEFEFEFEFEFEFEFEFEFEFE1B1A19405B40D2AD89121A40),
    .INIT_04(256'h65AEEE9D934A9B5BADF6129AA39B5BC989C9898989CA001AF5ECACECECEDF663),
    .INIT_05(256'h2323E32423E324242424246D6DB6F692D31C8BD4D3D4D4411C65F76E4A1C6565),
    .INIT_06(256'h1CD48B8BD41CD3D31CD425AEAEAED3D3ABECF4EC63A36363642323E323232324),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD3DC),
    .INIT_08(256'hFEFEFEFEFEFEF5B4F5F5FEFEFFFEFEFF24AD246DFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hA3ABECECABA3A3A3A3A362ABECECACACABA3A3ABF4FEFEFEFEFEFEFEFEFEFEFE),
    .INIT_0A(256'hADFEFE6463EDACA463636259A2EBABAAA3ACACB5FFFFF7EEF6F7F6B5F4F4F4F4),
    .INIT_0B(256'h005AC8404892B6FEFEFEFEFEFEF6FEFEFEFEFEF589ACA35AECC9AD64636440D2),
    .INIT_0C(256'h1CCA81C1020AA464F7AD12A3A35AC9C9C9898889C9898040EDF5A3A3F5F5F563),
    .INIT_0D(256'h2323232323242323232424242464641B1CD38BD4D3D4D34265AEF765421D2565),
    .INIT_0E(256'hD4D38BD31C1C8BD41CD3AEAEF75C8A64ECECF4AC63AC231B2323232423232323),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6ED31C),
    .INIT_10(256'hFEFEFEFEFEFEFEACB4F5FDFEFEFEFEAD24B6246DFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h63ABECACECA3A3A3A3A362ABECACABABABABF4F5FDFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_12(256'hFEFFB564EDA363ACACACACEBEBEBAB62ABACACFFFFF6A453E4F6FFFEF4F4F4F4),
    .INIT_13(256'hD21BA4ACF6FFFFFFFEFEFEFEFEF5FEFEFEFEFEF51BD11111126DADADADD1D263),
    .INIT_14(256'h1381D2135CEEF6ADF7645AA35AC989D2C989C9C98081C940D2F5F5ACECECF563),
    .INIT_15(256'h2323231BDADB232323DBDBDB242424242493D3D4D31C8A8B65AEF6258A651D6E),
    .INIT_16(256'hD48BD3D41DD48A1CDB65AEB7AED31BACF4F4F56C1B1B23232323242323232323),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDB1CD4),
    .INIT_18(256'hFEFEFEFEFEFEFEF5ACF5FEFEF5FEFE236DB56D6DFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h63ABECEBEBA2A2A2A2A262ABECECECF4F4F5F5F5F5F5FEFEFEFEFFFFFEFEFEFE),
    .INIT_1A(256'hD2F6F6ACA3A363ABECF4ECABA3ABABA3ABA3F6FFF6A4520009ADFFFFF5F4F4EC),
    .INIT_1B(256'hF6F6F6FEFEF6FEFEFEFEFEFEFEF5F5FEFEFEF6F6F56C1A0040B6FFF61AACF640),
    .INIT_1C(256'h5BA4EDEEF6AE6D64AD5B5B5AC9895B12C9C9C98081C989C940D1EDF5EDECF5F5),
    .INIT_1D(256'hDBDB23DBDADADBDBDB2324231B231BDB1C1CD3D3D3D4428B65AEB61CD3651C6E),
    .INIT_1E(256'h8BD3D31C1D8B931CDBAEAEAF65D264F4F5F5641B2323232424231B24232423DB),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6DD3D4D3),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_033792_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n60 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i33_008,inst_doa_i33_007,inst_doa_i33_006,inst_doa_i33_005,inst_doa_i33_004,inst_doa_i33_003,inst_doa_i33_002,inst_doa_i33_001,inst_doa_i33_000}));
  // address_offset=34816;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFF830FFDE7E1D3E08EFF1E6001FFFFFFFFE3FFFFEFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFF030F73C228FBF00EF0FEC000BFFFFFFFCDFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFF071FCF0036FFF81EB7FD80003FFF7FFF8FFFFFFFF001FFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFE171E00039FFFEC1EBFFB80001FFFFFFE0FFFE7FFF0003FFFFFFFFFFFF),
    .INIT_00(256'hFEFEFEFEFEFEFEFEF5F5F5ACF5F5FEAD6CB5FF6DB6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hA3ECECECECABA2A2A2A3A2A3ECF4F4F4F4F4F4F4F5FDFEFEFEFEFEFEFEFEFEFE),
    .INIT_02(256'hD2D2ADACA36263A3ABABABABACABA3A3A2ACF6F7A55349C052A4F6F6B5F5F4EC),
    .INIT_03(256'hF5F5F5F5F5F5F6F6FEFEFEFEFEFEFEFEFEFEFEFEF5FEFEF564F6FF6C63F663C9),
    .INIT_04(256'hA4EDE49BC180D265AE5B5BC9C9AD5CC9C9898081C9C989808988C9A3EDA3ECF5),
    .INIT_05(256'hDBDADB23231BDB1BDBE32323232323DBDBDBDBD31CD442D366AEB6D31C251C66),
    .INIT_06(256'h8BD31C1DDC8AD4D324AEAEAE1B1BB5F4AC1BDB24232423DBDB1B1B1B242423DB),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1CD4D38B),
    .INIT_08(256'hFEFEFEFEFEFEFEFEFEAC63ACF5F5FDFE6CB5FF6DB6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hA4ACACAC64631B6363636363ECF4ECACEBECF4F4F5FDFEFEFEFEFEFEFEFEFEFE),
    .INIT_0A(256'h5B11C9ACACA3A3A3ABABEBABABA3A3ABABADF6EE9C52099BEDF7FFF7F6EDF5AC),
    .INIT_0B(256'hECF4F4F4F5F5F6F6FEFEFEF6EDEDF5F6FEFEFEF6F5F5F5FEFEF6F6ADF56340D2),
    .INIT_0C(256'hD38180C04A9CADF6F65A1240AEAD40C9808089C9C989898189D2C98012C9A3F5),
    .INIT_0D(256'h23DBDBDB24231B2423DB232324232423DBDBDADBDBD342D4AEAEAED31C1C1D6E),
    .INIT_0E(256'hD3D41D1DD48ADCD36EB7AE65D3ADAD22D2DB24242423DB92DBDB1BDBDBDB23DB),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6EDCD48B8B),
    .INIT_10(256'hFEFEFEFEFEFEFEFEFEF5ABECF4F5FDFEADF6FF6D6DFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h92DBD3D392939393DBD3DB1A63ACF4F4F4ECF4F4F5F5FEFEFEFEFEFEFEFEFEFE),
    .INIT_12(256'h515B1B1AEDABA3A3ECECABEBABA3A3631B64F6EEA452A4EEF7F7F7F6F6F6F563),
    .INIT_13(256'hECF4F5F5F5F6FEFEFEFEFEACC04909F5FEFEFEFEF6F5F5F5FEFEFEAD630089C9),
    .INIT_14(256'hD31465A5ADADADB6F51A40ADFFD240C1C9C9C98988898989CACAC9C9804012ED),
    .INIT_15(256'hDB2323DB2324241B24241B242424232423DADAD2D3924A1CAEAEAE9365DC25AE),
    .INIT_16(256'hD41C1D1C8BD3D31CAFAE651C1C64D2D223242424DB928992DADADBDBDADB2423),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1CD4D38AD3),
    .INIT_18(256'hFEFEFEFEFEFEFEFEFEFEF4ABF4B4F5FEF6FEFFB66DFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h9B939C949494949CDCDCDBD3D3DA1B64ACF5F5F5F5F5FDFEFEFEFEFEFEFEFEFE),
    .INIT_1A(256'h115AAD1B1BEDA3ABEBABA3ABA3631A92DC65F6F6A463EDF6EEEDEDA4A4F6F6AE),
    .INIT_1B(256'hF5F5F5F5FEFEFEFEFEFEFEA392D251F6FEFEF6F6F6F6F5F5F6FFADC9408989C9),
    .INIT_1C(256'h65B6AE6D242CB5FEF6C91BFFAD40C9CACAC989898989C9CACA8989898989405B),
    .INIT_1D(256'h241B232324246D242324241B24242CDB242392DBD3D3411CAEAEAE9365D365AE),
    .INIT_1E(256'hDC1D1C1C8AD38B66B76E1CDB9292D2DBDBDBD2499192DADADBE3232323DBDB24),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAED4D38B8A1C),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_034816_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n60 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i34_008,inst_doa_i34_007,inst_doa_i34_006,inst_doa_i34_005,inst_doa_i34_004,inst_doa_i34_003,inst_doa_i34_002,inst_doa_i34_001,inst_doa_i34_000}));
  // address_offset=35840;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFE1E3E0043DFFF761EBFFB80000FFFFFFC0F7F9BFFF80787FFFFFFFFFFF),
    .INITP_01(256'hFFFFFFC3E3809FBFFFF7B1FBFFB308017FFFFFC0FFF31FF780A807FFFFFFFFFF),
    .INITP_02(256'hFFFFFFC3E043FFFBFFFBD9FBFFF700073FFFFF86FFE60FFF83F801FFFFFFFFFF),
    .INITP_03(256'hFFFFFF83C013FFFDFDFDCDFBFFFE001E3FFFFE06FF8407FF9F07007FFFFFFFFF),
    .INIT_00(256'hFEFEFEFEFEFEFEFEFEFEFEB4F5F5FDFEFEF6FFB66DFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h254A9394DCDCDCDDDD251D1D1DDCDC93DB1B64ACF5F5FDFDFEFEFEFFFEFEFEFE),
    .INIT_02(256'h1212ADF6D2ACECABECA3A3AC1B8A932525DC6DF6ACADEEAD5B5B530A09A4F6FF),
    .INIT_03(256'h5BF5F5F5F6FEFEFEF6FEFEAC5A92E4FEFEFEFEFEFEFEFEFEFFFED24089898181),
    .INIT_04(256'h5B64236CB5FEFEFFFE89ADFF1280C981C981808081C9CACAC989898989894000),
    .INIT_05(256'h6D2423242424646D24246C1BDB246C24DB6C23D2DBD34924AEAE6DD365D365AE),
    .INIT_06(256'h1C251CD48AD31CAEAE241B92499192DADBDBDADADA23DBDBDBE323232324DB24),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF65D38B8AD31C),
    .INIT_08(256'hFEFEFEFEFEFEFEFEFEFEFEFEB4F5FEFEFEF6FFB66CFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hAE8AD4DCDCDCDCDC1DDC1DDD1DDDDDDDDCD3928ADB6CB5FEFEFEFEFEFEFEFEFE),
    .INIT_0A(256'h111A64F6AC1AF5ACABA3A31B8ADC2525DC4A9265ADEDEEA452090901C05BF6FF),
    .INIT_0B(256'h8A1BEDF5F5F5FEFEFEFEFEF5A4EDF6FEFEFEFEFEFEFEFEFFFE1B40C980C9C981),
    .INIT_0C(256'h1AACF5FEFEFEFEFEFEDAF6F64080121B894089C90ACAC98988C9C9C98040DB24),
    .INIT_0D(256'h246D24242324246C6D242464DB1B246C24926C23D2DB8A25AEAE651C25D36EAE),
    .INIT_0E(256'h1D251CD393931CAE65DBDB89DA92DBDB23DBDB232323232323DB242423232423),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7D3938B8A1C1D),
    .INIT_10(256'hFEFEFEFEFEFEFEFEFEFEFEFEF5ACACF4FEFEFEB66CFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hAE8A8A93D4DC1D251D1D251D1DDDDDDDDDDDDDDC938AD364F6FEFEFEFEFEFEFE),
    .INIT_12(256'h095A64EDF51A6CF5AC631B93DD2525DC934A4A001BEDED9C52524A4A099BEDF6),
    .INIT_13(256'h92405BECF5F5FEF6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFFF61240C98940125B89),
    .INIT_14(256'hACFEFEFEFEFEFEFEFE64FFAD0064F76480D2D1D2C9C9C9C9C9898040891C6E6E),
    .INIT_15(256'h246C6D23242324246C6D242424DA23246C2392641BDB9265AEAE651C1DD4AEAE),
    .INIT_16(256'h651D1C939392D3DBD22392DBDBDA2324231B2323242323232424246C24DB2324),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF658B8B8A8A1D1D),
    .INIT_18(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEACABA36CFEFEAD6CFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h6E93DC1D25252525DDDDDDDDDD1D1D1CDCDDDDDDDDDDDDDCDCADFEFEFEFEFEFE),
    .INIT_1A(256'h115AA4ECACAC1BF5ACDA93E5E51DDB938A4A4A0092ADED9B53525253EDA4A4F6),
    .INIT_1B(256'h0A411B63ECF5F5FEFEFEFEFEF6FEFEFEFEF6FEFEFEFE644080C9C988805BAD89),
    .INIT_1C(256'h75FFFEFEFEFFFFFFFFB5FE2424FFAE40C08080888080808080C9D21B656E6E9C),
    .INIT_1D(256'h64246D242324DB24246C6D2424249223246DDB92241B9224AEAE651C1CDCAEAE),
    .INIT_1E(256'h651DD48B8A929291DBDBDB23DADB23232424242424242424242424646424D223),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7DC938A8A8B651D),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_035840_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n60 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i35_008,inst_doa_i35_007,inst_doa_i35_006,inst_doa_i35_005,inst_doa_i35_004,inst_doa_i35_003,inst_doa_i35_002,inst_doa_i35_001,inst_doa_i35_000}));
  // address_offset=36864;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFF83C0A7FFFCF6FCE4FFFFFC01FE1FFFF806FF8807FFBC80003FFFFFFFFF),
    .INITP_01(256'hFFFFFF8380EFFFFE7A7E727FFFFDFFFE07FFE00EFF9003FF8100001FFFFFFFFF),
    .INITP_02(256'hFFFFFF0781EFFFDC393C307FFFFFBFFE01FFC4FEFF9003FF00000027FFFFFFFF),
    .INITP_03(256'hFFFFFF0781EFFF6E1C0E187FFFFFFFFE003C77FEFFA001FC0201001BFFFFFFFF),
    .INIT_00(256'hFEFEFEFEFEFEFEFFFEFEFEFEFFFEB5F563ACFE6C24FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h25D41D252525DCDC1DDC9393DCDCDDDDDDDDDDDDDDDDDDDDDDDC25F6FFFEFEFE),
    .INIT_02(256'h115AA4ACACEC63AD2593DDDC1CDC94934A4A4A414964ADA45B52529BE5A4A4F6),
    .INIT_03(256'h4A0A4A1B5BA3F4F5FEFEFEFEFEFEFEFEFEFEFEFEAD920089CAC9898980A4F540),
    .INIT_04(256'hADFEFEFEFEFEFEFEFEFEFE6CFEFF9200DADB0000408ADB24656E6E256E6E2500),
    .INIT_05(256'h24646C6CE32424DB23236D6D2424DB91236C6C92D224DADB65AE25251C1CAEAE),
    .INIT_06(256'h661CDB8A9292929224DB24DBDB2424242424242424242424232464246C24DB92),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAE8BCB8A8AD3651D),
    .INIT_08(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFDB4FD6BFDFE6CFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h25DCDCDCDCDCDC1DDC93494A938B94DCDDDDDDDDDDDDDDDDDDDDDC1CB6FFFEFE),
    .INIT_0A(256'h125BACACA3ECAC6424DCDC1CDC93DC4A9293494A00DBADADA49B5B9B5B64F6EE),
    .INIT_0B(256'h0A4A0A41D31B63EDF5FEFEFEFEFEFEFEFEF66CD20040CAD289C9C9C912F6F640),
    .INIT_0C(256'hADFEFEFEFEFEFEFEFEFEFEB6FFB6DBAEFEAD1B65AEB6B7B7B6B66E6E6E6E6D49),
    .INIT_0D(256'hD3236C6D24DA24DBDB23246D6C2323DA92236C2392DB23D2DBAE25251C1DAEAE),
    .INIT_0E(256'h66D4D38A929292DB241B24DB24242424246C242424242424242323646C242392),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF258BD38B8ADC6565),
    .INIT_10(256'hFEFEFEFFFEFEFEFEFEFEFEFEFEFEFEB5F5FDB5FEB6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hDCDCDCDCDCDDDDDCDC49014A93DCDDDCDCDCDDDDDDDDDDDDDDDD1DDCDC6DFFFE),
    .INIT_12(256'h1263EDABA3ECAD2425D4DC2593DC934ADB4A4949410064F6F6EDA5A5A5EEAE1C),
    .INIT_13(256'h014A4A4A0193D31BA4F5FDFEFEF6F6AD65654000C909C0801B5B1212A4FFAD80),
    .INIT_14(256'hADFEFEFEFEFEFEFEFEFEFFF7FF64A5F7AD81A4FFFFFFB7B6B6B6AE6E6E6E6E8A),
    .INIT_15(256'h49DB236C6DDADA23DBDB23246C24DBDB91922464DBDBDBDB926D1C1D1D25AEAE),
    .INIT_16(256'h66D3D38A92929224232424DB6C242464246C246C232464642324DB246C6CDBDB),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD3D3D38A8A1C6565),
    .INIT_18(256'hFEFEFFFFFFFEFEFEFEFEFEFEFEFEFEFEB5FEB5FEFEFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h9393DCDCDDDD25DC4A019394DDDDDD1DDD9493DCDCDCDCDDDDDDDD1D1DDC6DFE),
    .INIT_1A(256'h5BEDEDA3A3AC6C2525932593DCDC01DCDB0149494901411CADEEEEAEAD65DB41),
    .INIT_1B(256'h014A4A4A4B0A4AD3D2DB246D6D24DCDCDBAEB66481125BADED1A12A4FFFF6480),
    .INIT_1C(256'hACFEFEFEFDFEFEFEFEFFFFF7B6AD1B5BE5E5125CF6FFFFF7B6B6B6AE6E6E6E93),
    .INIT_1D(256'h9292DA246D2449DBDBDBDBDB246C1BDBDA49DA6C23DBDBDBD26D241D1D65AEAE),
    .INIT_1E(256'h65D3938A9292D224236424DB6D24246C246C6C6C1B246C6CDB6C23DA246D1BDB),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF793D3D38A8A1C656E),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_036864_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n68 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i36_008,inst_doa_i36_007,inst_doa_i36_006,inst_doa_i36_005,inst_doa_i36_004,inst_doa_i36_003,inst_doa_i36_002,inst_doa_i36_001,inst_doa_i36_000}));
  // address_offset=37888;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFF0781FFFF660C460A7FFFFFFFFE00027FFCFF480070041B0005FFFFFFFF),
    .INITP_01(256'hFFFFFF0381DFF7B60C02025FFFFFFFFF00007FFDFB4000000C360002FFFFFFFF),
    .INITP_02(256'hFFFFFF8383FFF7B20623031FFFFFFBFF00007FFFF8920000186C0C017FFFFFFF),
    .INITP_03(256'hFFFFFF8383FBF7980601011FFFFFEDFF80027FFFF082000030DC2C001FFFFFFF),
    .INIT_00(256'hF6F6F6F6FEFEFEFEFEFEFEFEFEFEFEFEF5F5F5F5FEFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h93DCDCDCDC25DD934A8BDC1D1DDD251DDC93934A93DCDCDDDDDDDDDDDD1DDC25),
    .INIT_02(256'hACF6ACA3AB632425DC1DDC931C934ADD924A4949014949008A1B241CDB4A8A8A),
    .INIT_03(256'h014A4A4A4A4B4B4A4B0A0A5394DC25DD936DB6FFAD64F6F65B5BEDFFFFF6C981),
    .INIT_04(256'hACFEFDFEFEFEFEFEFFFF6E6E6EF6F6A553A5ED5B53F7FFBFBFB6B6B66EAEB6DC),
    .INIT_05(256'hDB4992DA6C6C9192DB1BDBDBDB2424DADB9289DB24DB24D292641C1D1C65AEAE),
    .INIT_06(256'h658A92899292DB24246C23246D24246C246C6C641B646C6DDB236CDBDA6C2492),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF793D3D38A8A1C65AE),
    .INIT_08(256'h1CAEF6F6FFFFFFFEFEFEFEFEFEFEFEFEFEF5F5F5F6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hDCDCDCDC2525934A4BDC1D1DDD2625DC94D49393DCDDDDD4DDDDDCDCDDDD1DDC),
    .INIT_0A(256'hF5F4A3A363DB2525DC2593DCDC01DCDD4A4A4949010149490001418A934A4A93),
    .INIT_0B(256'h014B0A4A4A4B4B4B4B549C9DE5E6DD4BDC6E6DFFFFFFB624ACFEFFFFFF6380AD),
    .INIT_0C(256'hACF5F5FDFEFEFEFFF66D25251D25AEF7F65C64EE535BF7FFFFF7B7B6B6AEB725),
    .INIT_0D(256'hD2919192236DDA49DADBDB9ADBDB24DAD2D24992DBDB24DB921BDB1D1C65AEAD),
    .INIT_0E(256'h654A92499292DB24246CDB246C236464246C6C64DB646C6D1BD26D2491236C91),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD4D3D38A8BD465AE),
    .INIT_10(256'hDC1CA4EDFFFFFFF6FEFEFEFEFEFEFEFEFFFEB4F5FEFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h93DCDC2526D44A93DC2525DC2525DCDCDC9393DC1D25DDDDD494DCDCDDDDDD1D),
    .INIT_12(256'h6BACABA31BD3DCDC25D49325934A25DC494A4901414901494A4A8A9293939394),
    .INIT_13(256'h4A4A524A4A4B4B0B0B5394DDDD9C94DDDC6E6EFFFFFFFFF6F6FFFFFFB523FEFE),
    .INIT_14(256'hACF5F5F5F6FEFEB66D25252525251C65B5F6125CE681A4FFFFFFB7B6B6B6B7B6),
    .INIT_15(256'h89DA9192DA6C234992DA23DADAD2232392DB924992DB232492D2931C1C65AE6D),
    .INIT_16(256'h6549929192922324236C1B246C236C24236C6C24D2646C6C2391246DDA9224DA),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1C8BD48B8BD465AE),
    .INIT_18(256'hDDD48A13A4EDEEF6FEFEFEFEFEFEFEFEFFFEF5F5FEFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hDCDC256EDC9393DC1D25DC256E1DDCDD939325DC2625DDDCDCDB4AD4DCDDDDDD),
    .INIT_1A(256'h6BABAB63D2938ADC254BDCDC4ADC2594494A414149414149494A4A924A939393),
    .INIT_1B(256'h1D0153534B4A4B534B94DCDC94DC25DC9325B6FFFFFFFFFFFFBEBEFFB6FFFEFD),
    .INIT_1C(256'hABF5F5F6FEFEB665652525252424641B2264A581A5A4C1F7FFFFFFB7B7B6B7F7),
    .INIT_1D(256'h40DA9291912464929192DBDB9292DB23929292499292DB24DB92D21C1C65AE65),
    .INIT_1E(256'h65494992929223241B641B246CDB24241B6C6C2492246D6C2392926D2389DBDB),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6E41D4D38BD465AE),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_037888_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n68 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i37_008,inst_doa_i37_007,inst_doa_i37_006,inst_doa_i37_005,inst_doa_i37_004,inst_doa_i37_003,inst_doa_i37_002,inst_doa_i37_001,inst_doa_i37_000}));
  // address_offset=38912;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFF83837B77980211019FFFFFF7FF80047FFFF1260000219A5880CFFFFFFF),
    .INITP_01(256'hFFFFFFD3035B73882110009FFFFFFEFF80007FFFE12600006334190087FFFFFF),
    .INITP_02(256'hFFFFFFD3835873083180008FFFFFFFFFC0007FFFE2460000C370B21007FFFFFF),
    .INITP_03(256'hFFFFFFC383403300318000DFFFFFFF7FC0007FFFE4440001C279360003FFFFFF),
    .INIT_00(256'h1D1DDCCA0A09A5F7F6FEF5FEFEFEFEFEFFFEFDF5FEFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hDCDC6EDC9393DD1D25DCDC6E25DC1DD44A25DC2526DDDCDD259393D4DCDDDDDD),
    .INIT_02(256'hABABAC1A92939325D39325934A2525934A49494141414949494A4A4A93938BDC),
    .INIT_03(256'h6F01534B53530A53949C9C9CDD26E54A5325FFFFFFFFFFFFFFFFFFF6FFFFFEFE),
    .INIT_04(256'hABF5F5FEF7AE6D6566656524636463A3A363AD6481E552A5FFFFFFFFFFB7B6FF),
    .INIT_05(256'h4991914949921BD29191DB239292921BDA91DA49929292232391D31C1C65AE65),
    .INIT_06(256'h1C49899292922324DB641B2424DB2424DB6C6C2489236D2C24924924249192DA),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB74AD4D48BD3656D),
    .INIT_08(256'h1DDDDDD4CA9CEDF6F6FEFEFEFEFEFEFEFFFEFEF5FEFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hDC2525DC93DC1D25DCDC2566DC1DDC4ADDDDDC2525DCDD2694DCDDDCDC8BDDDD),
    .INIT_0A(256'hACAC648A934ADC2493DC254B9325254A4A49494149494149494A4A93938ADCDC),
    .INIT_0B(256'hFFDC01945353534A4A4B5394DDDD944A0A6EFFFFFFFFFFFFFFFFFFFFFFF6FEFF),
    .INIT_0C(256'hACF5F6F66E6E6E6E666564ACACACABABECEC6CAE139CE5CAF6FFFFFFFFFFB7B7),
    .INIT_0D(256'h499163D24992DB1B91499223D29292DBDB919292499291DB2492D21C1C6EAE65),
    .INIT_0E(256'hD349499292922324DB6DDB2424DB232492246C2491DA6D24239249DA24929292),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1C8A1D8BD32565),
    .INIT_10(256'hDDDDDCD4935CEEEDF6FFFFFFFEFEFEFEFFFEFEF6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h2525DC93DCDC25259325661DDDDD4ADC25942525DCDC66DD93DDDD1D934A94DD),
    .INIT_12(256'hF5ED1B8A929325DC9325DC4ADC651D4A4A494901494949494A4A93924ADCDC93),
    .INIT_13(256'hFF6E024B949C9C9C934A539CDD94534B0176FFFFFFFFFFFFFFFFFFFFFFFFA4A4),
    .INIT_14(256'hB5F6B6AEAE6E6E6E6E6564ACACACECF4F5F5B5ADAD13ED5B64FFFFFFFFFFFFB7),
    .INIT_15(256'h4989641B0092DB6C1A8949DBD2899292DB899292499291DA24DB92DB25AFF7AE),
    .INIT_16(256'h24924992919224239264DB2323DADBDB92246D2391496D6CDB92498924DA8992),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAE411D8BD31C65),
    .INIT_18(256'hDDDDDCDCDC9313125BF6FFFFFEFEFEFFFEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h2525DCDCDCDC2593DC2625251D938B25D4DC2525DC25254ADCDDDDDD93DDDCDC),
    .INIT_1A(256'hA46425DC491CDD94DC259393DC6EDC4A49494901494949494A93924ADCDC9325),
    .INIT_1B(256'hFFFFDC024B539C9CDCDCDCDDDD94940BDBFFFFFFFFFFFFFFFFFFFFFFFFAD12E5),
    .INIT_1C(256'h6D6D6E6E6E6E6E6E6D64ACF4F5F5F5F5F5ECF5F5B6655CE5C1EEFFFFFFFFFFFF),
    .INIT_1D(256'h5248A4A40052D2AD1BD289DBDB499192DB919192499291912323DB246E6EAEAE),
    .INIT_1E(256'hAED349929192231B9264DBDBDB9292DB92DB6C239200246DDB924949DBDB4991),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD3D4D48B1C1C),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_038912_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n68 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i38_008,inst_doa_i38_007,inst_doa_i38_006,inst_doa_i38_005,inst_doa_i38_004,inst_doa_i38_003,inst_doa_i38_002,inst_doa_i38_001,inst_doa_i38_000}));
  // address_offset=39936;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFEB814031003180007FFFFFFFFFE000FFFB644C000184F26CA000FFFFFF),
    .INITP_01(256'hFFFFFFE9C00031803180007FFFFFFFFFE000FFF6E48C000388E278600CFFFFFF),
    .INITP_02(256'hFFFFFFF1C000101281E0007FFFFFFFDFF001FFFDE88C000308C478C0007FFFFF),
    .INITP_03(256'hFFFFFFF4C00010120060007FFFFFFFEFF001FFBBF00C0006018470C0007FFFFF),
    .INIT_00(256'hDDDDDDDDDDDDD3D25BA4EEF6F6F6FEFEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h25DCDCDCDC25DC932526251DD3011DDC932525DD252693931DDD25DDDCDDDCDC),
    .INIT_02(256'hC9AEB7DC9325DC93DC1C9393256E934A494909014949494A924A01DCDC93DC25),
    .INIT_03(256'hFFFF6E01544B0A53949C9C9C9C9CDD0A6EFFFFFFFFFFFFFFFFFFFFF7A5C1EDED),
    .INIT_04(256'h25252525252525252464F5F5F5F5F5F5F4F5F5FEB5F664E59C12FFFFFFFFFFFF),
    .INIT_05(256'h9289ACAD8949DBF664D292DADB899149D291499249929249DB24246D65252525),
    .INIT_06(256'hAEDB00929292DB1B4924DBDBDB9292D2919124239248DB64DB928989D2DA9189),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF65D31C8B1C1C),
    .INIT_08(256'hDCDDDDDD1D1DDCD35B5B5BA5EDF5FEFEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h1CDCDCDC1DDC4ADC252525DC01D3254ADC25251D66DC42DCDC2525DCDC4A4AD4),
    .INIT_0A(256'hADFFB693DC25DC9325DC93932525934A494A49014949494A4A01D4DC93DC2525),
    .INIT_0B(256'hFFFFFFDC4B9C949494949C9DE5E69CDCFFFFFFFFFFFFFFFFFFFFF75CC1E5E480),
    .INIT_0C(256'h252526252566656564B5F5F5F5FDFDB5ACF5FEFEFEF6F65CE50A64FFFFFFFFFF),
    .INIT_0D(256'h92D2ACADD200DBF6ACD2DAD2D2919149929249924989924992246D6E25252525),
    .INIT_0E(256'hAE2400929191DBDB49DBDB92DB92928991491B23929192231B9191D2D2D2DA89),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB68A1CD3D31C),
    .INIT_10(256'hDCDDDDDDDDDDDCD3D25B52A4F6F6FEFEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hDCDC93DC1D934ADD2625DC4A4A25D392DC252525254A93DC1D25DDDC93004AD3),
    .INIT_12(256'hF6AD659324DC93DC25D48BDC2525934A494A494149494A4A0193D48BDCDC2525),
    .INIT_13(256'hFFFFFF6E01939CDDDDDDE6E6E5E5536FFFFFFFFFFFFFFFFFFFF71B13E59C8064),
    .INIT_14(256'h252525656D6E6524ADFDFDFEFDFEF5ACF5FEFEFEFEF6F6AD53A5C1EDFFFFFFFF),
    .INIT_15(256'h1BD2DADB8948D26C641A1B92929292499291499249899249916CAE6E25252525),
    .INIT_16(256'h6D2400929192DBDB4992DB92DB9249499289D2239291D2DBDB919264D2D26489),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1CD4D48B1C),
    .INIT_18(256'hDDDDDDDDDDDDDC93CA1B63EDF6F6FEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hDC93DCDCDC4A932566DC9301D31C4AD3DC252525D349DCDC251DDCDB00494A93),
    .INIT_1A(256'h6464641CDDDC93DCDC9493DC6625524A4A4A4141494A49494A934AD4DC2526DC),
    .INIT_1B(256'hFFFFFFFF9C4A549494DDDDDDDD93DCFFFFFFFFFFFFFFFFFFEED29CEE9C81A5F6),
    .INIT_1C(256'h2525666D6D6E6524F6FDFDFDFEFEF5F5F5FEFEFEFEFEF6F71B5CE5C1ADFFFFFF),
    .INIT_1D(256'hD249000000490040D21B6392899292089149499249929289916DAE6525252525),
    .INIT_1E(256'h65240089919192DB89919291929249929189DA23DA92D2D2DB9192ADDAD2B5D1),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAED31D8BD3),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_039936_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n68 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i39_008,inst_doa_i39_007,inst_doa_i39_006,inst_doa_i39_005,inst_doa_i39_004,inst_doa_i39_003,inst_doa_i39_002,inst_doa_i39_001,inst_doa_i39_000}));
  // address_offset=40960;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFF4C000101E0020007FFFFFFFBFF803FF77F90800060180E080203FFFFF),
    .INITP_01(256'hFFFFFFFEC000583FC000087FFFFFFFDFFC07FFFFF908000C0300C100003FFFFF),
    .INITP_02(256'hFFFFFFFEC0076CBFC0000CFFFFFFFFFFFC07FFFFF808001802008160001FFFFF),
    .INITP_03(256'hFFFFFFFF60038EFFC0800CFFFFFFFFFFFE0FFFFFF818001800018278000FFFFF),
    .INIT_00(256'hDDDD1DDD94935252538A64F6FEF6FEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h939CDDDC9200DC661D8B4A01DC934ADC1D251DDC8A93DCDD25DCDC4A01494993),
    .INIT_02(256'hACF5AC6D1CDC9325DC9393DC66DC934A494941494A09494A934A93DCDD2625DC),
    .INIT_03(256'hFFFFFFFF6E0A939494949CDD9C4AB7FFFFFFFFFFFFFFF7A4C9A5EE9BC1EDF66D),
    .INIT_04(256'h256E6E6E6E6E24B5FEFEFDFEFEF5B4F5F6FEFEFEFEFEFEF6EE81A4ED0AA5FFFF),
    .INIT_05(256'h489200494949490000931C8949DA92419249498949919249926D6D6525252525),
    .INIT_06(256'h65654949919291DB9249929292929189DA898964DB91D2DB9292D2ED1A23B589),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDC1CD3D3),
    .INIT_08(256'hDCDC934A4A4A4A9393931BEDF5F6FEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h93DCDC9B4A4A2525934A0192DC4993DC2525DC939293DC25DCDCD3004A494A93),
    .INIT_0A(256'hFEF5B56D24D4DC25DC9393DC6EDC934A4A494149490109934A4ADCDC2525DC93),
    .INIT_0B(256'hFFFFFFFFFF25DD9D9CDDDD9C0125FFFFFFFFFFFFFFAD125BEEEE5313F6F7ADB5),
    .INIT_0C(256'h6E6EAEB7AE6D6DFEFEFDFDFEFEF5F5FDFEFEFEFEFEFEFEFEF6A581A5EE9C13AE),
    .INIT_0D(256'h6D1B4900494848494900899248DB9200498940DA6D899292DB6D6D6565652566),
    .INIT_0E(256'h25659248919249DA9249919292DBD289D21B001B6CD1D1DBDB4812F5636CF61A),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6E1C1C8B),
    .INIT_10(256'h934A0149494A939393DC931CADFEFEFEB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hDCDCD392019325934A4A01939349D3DC66DC93939392DC25DC1C1BC940414A93),
    .INIT_12(256'hFEFDFEAD2593DCDDDC9393DC65DC934A4A49494949494A924A93DC2526DCD34A),
    .INIT_13(256'h1BADFFFFFF76DDE5DDDD9D4B93B7FFFFFFFEF6A51313ADEEE5019CFFFFF6FEFE),
    .INIT_14(256'h6EB6B7B7B665B5FEF5F5FEFEF5F5F6FEFEFEFEFEFEFEFEFEF5ADAD125BEEED12),
    .INIT_15(256'hB66DD300494849000000404849DB9241499289DBF61B0092246E6D6565656E6E),
    .INIT_16(256'h1C65DB0049924992D2494949891B1B1A88231B89ACACD2D223891AF5ACADF663),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1C65D3),
    .INIT_18(256'h49014949494A9393DCDC9393B6FEFEFEB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hDCD4934A00DCDC4A4A4949924A93931D65D35293934A25DDDC1B63A31B894A92),
    .INIT_1A(256'hFEFEFEB56593DDDD944B93252593934A4A4941014A4A4A4A93DCDC661D939393),
    .INIT_1B(256'hE4531BA5FFFF25DDE5DDDD9465F6AE645B13129CE5EEED530AEDFFFEB6FEFEFE),
    .INIT_1C(256'hB6B6B6B66D6DFEFDF4FDFEFDF5F6FEFEFEFEFEFEFEFEFEFEFE6CADEEA412A5EE),
    .INIT_1D(256'hFEF6DC004948494924D3DB9192DB494949DB92D2F66400DB6D6E6E6E6E6E6EAE),
    .INIT_1E(256'hD3652449499249499291494948D21B636391DB891AF5B5D21A1A1AF5ACF5F6AC),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF651C1C),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_040960_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n76 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i40_008,inst_doa_i40_007,inst_doa_i40_006,inst_doa_i40_005,inst_doa_i40_004,inst_doa_i40_003,inst_doa_i40_002,inst_doa_i40_001,inst_doa_i40_000}));
  // address_offset=41984;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFD600387FFE0E04DFFFFFFFFFFF70FFFFFFA180030000102FC000DFFFF),
    .INITP_01(256'hFFFFFFFFB00183FFECF00DFFFFFFFFFFFE1FFFFFFA180060000000FE0081FFFF),
    .INITP_02(256'hFFFFFFFEB80603FFFDB009FDFFFFFFFFFF19FFFFFE100040000001FF80803FFF),
    .INITP_03(256'hFFFFFFFFD80307FFFFA02008FFFFFFFFFB3FFFFFFE100080000001FFC0841FFF),
    .INIT_00(256'h4A4A4901014A9393DCDCD4DC1C1CDBB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hD4938A4941DC934A4A494A8A4A939325DC934ADC4A9225DC1C63A3A3A35B8949),
    .INIT_02(256'hFEFEFEF665DC25DD934B932525939349494101494A4A4A4A93DC252593934ADC),
    .INIT_03(256'hA4EDE55BC9A56525E5E5DD8B1C645CA5EEEEEEEEE5530AA4F7FFB6F6FEFEFEFE),
    .INIT_04(256'hADADADB6ADF5F5F4F5FEFEF5FDFEFEFEFEFEFEFEFEFEFEFEFEF56CACF6F65C5B),
    .INIT_05(256'hFEFF6D0089914949F7FF6DDB4992494949239189F66C00246E6E6E6E6E6E6EAE),
    .INIT_06(256'hD31D65D30092924991924992924063631B4900000064FEF5636323F5F5F6F6F5),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7DC65),
    .INIT_08(256'hCA8A4949418A92931DDCDCDDDDDC8A6DFFB7B7FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h934B4A014A934A4A928A8A49929293E5934993DC0093DCDC1C5BA3ECECAC63D2),
    .INIT_0A(256'hFEFEFEFE65DC1DDD934A93252593934901494949494A4A93931D2593934A93D4),
    .INIT_0B(256'h64139CEDA55313DCE5DDDC5CEEEEA5ADA5A55B1213A4F6FFF6ADFEFEFEFDFEFE),
    .INIT_0C(256'hB5B5F5F6F5F5F5F5FEFEFDF5FEFEFEFEFEFEFEFEFEF5FEFFFEFDF4F5ACF5F6ED),
    .INIT_0D(256'hFEFFB6406C1A0000B5F66D230092494992DB9291B56489646D6D6D6E6D6D6DAD),
    .INIT_0E(256'h1CD46E654949924949928989DBD288AC1B0048490092B5FEF5AD6CB5F6FEFEFE),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2524),
    .INIT_10(256'h5BD39249498A4AD425DCDCDDDDDDD4934A8A24B7FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h8B4A49494A4A01499289924AD38ADCDC8A01DCDC0093941C5BACECECECECECA4),
    .INIT_12(256'hFEFEFEFE251D1DDC934A9325DDD392010149490149494A93D425DC934A4A9393),
    .INIT_13(256'hF7F6A41B135CA51CDC938A5B53CAD31B5C64ADF6F6FEF6ACADFEFEFEFEFDFEFE),
    .INIT_14(256'hACACADF5F5F5ACFEFEFEFEFEFEFEFEFEFEFEFEFDFDF5FEFFFEFEF5FDFEF5B5F5),
    .INIT_15(256'hFEFEFE23F66C001AADDA6C230092494992DBDBDA64DBD2246525256D6D24DB24),
    .INIT_16(256'h65D365AE1C00924949499249921B1AD2920040490000B5FEFEFEF6F5FEFEFEFE),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6DB),
    .INIT_18(256'hA45BD20049924ADC25DCE5DDDD1DDCDCDC93DC6EFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h8B4989924A4A49D2898A92008A8AD393498ADC930093942464EDF5F5F4F4ECEC),
    .INIT_1A(256'hFEFEFEFE6D1D25DC934AD325DDD44A0149494941494992931DDD939301939393),
    .INIT_1B(256'hB6F6F6F6A5D35C1C8A4264EDEDAEF6F6FEFFFFFEF6ADACF5FEFEFEFEB5FEFEFD),
    .INIT_1C(256'h63ACB5F4F4ACF5FEFEFEFEFEFEFEFEFEFEFEFEFEACF5FEFEFEFEF5FDFEFEFEF6),
    .INIT_1D(256'hFEFEFFAD23F5B4FEAC00B5DB00924991DADB24DADB4992DBDBDB92DB24DA91DA),
    .INIT_1E(256'h651CDC6E658A4A8A4949929249D2646489004000DB6DB6FEFEFEFEFEFEFEFEFE),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF24),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_041984_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n76 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i41_008,inst_doa_i41_007,inst_doa_i41_006,inst_doa_i41_005,inst_doa_i41_004,inst_doa_i41_003,inst_doa_i41_002,inst_doa_i41_001,inst_doa_i41_000}));
  // address_offset=43008;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFDC01C7FFF3A06008FFFFFFFFFF7FFFFFFE100080016001FFE1A49FFF),
    .INITP_01(256'hFFFFFFFFFC00E3FFF8006008FFFFFFFFFFFFFFFFFE100000236001FFF1AC8FFF),
    .INITP_02(256'hFFFFFFFFEC00EFFFFFE0E00CFFFFFFFFFFFFFFFFFE10000023F081FFF13CCFFF),
    .INITP_03(256'hFFFFFFFFFE00FDFFFFE0E00CFFFFFFFFFFFFFFFFFE30000027F081FFE33CCFFF),
    .INIT_00(256'hE3A35BD24952931D1DDC25DDDD1DDCDC25949325FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h4A00D2924A09D25B89641B9192494A4A40DBDC4A4192DC1CADF5F5F5F5F4F4EC),
    .INIT_02(256'hFEFEFEFE6D2525948B4ADC25DCDC49494A494949494A8ADC1D93934A4A939393),
    .INIT_03(256'hFFFEF5F6F6AD641C8A6EFFF6B6B6F6FEF6F6FEF6F5F6FEFEFEFEFEF5F5FEFEFE),
    .INIT_04(256'h63B5B5F4ACACFEFEFEFEFEFEFEFEFEFEFEFEFEFDABFEFEFEFEFEFDFEFEFEFEFF),
    .INIT_05(256'hFEFEFFAD00DAAC6C23D2ADDB00929192DB2424DB92499292929292DB24DB91DA),
    .INIT_06(256'h1C65D365AE1C0192924992494949916CAC234900DAB5B5FEFEFEFEFEFEFEFEFE),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6),
    .INIT_08(256'hECA3A35B494A93251DDC25DD1D1DDCDC25DC93DCB6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h4A001BD209001B1AD2AD1BDAD34A92494892DC4A4992DC1CEDF5F5F5F5F5F5F5),
    .INIT_0A(256'hFEFEFEFE6D2525948A4ADC25DC93014A4A494949498A93DC939393019293934A),
    .INIT_0B(256'hFEFEFEFEF6ADADAD64AEADB5F6FEFEFEFEFEFEFEFEFEFEFEFEFEFEF5FEFEFEFE),
    .INIT_0C(256'h23ADF4ACACFEFEFEFEFEFEFEFEFEFEFEFEFEFEACABF5FEFEFEFEFEFDFEFEFEFF),
    .INIT_0D(256'hFEFEFEB51B91894889D2DBD341929289DB6424DBDB4992929292929224DB91D2),
    .INIT_0E(256'h24651C1C6E658A8ADB9249524949899163F51B48894023FEFEFEFEFEFEFEFEFE),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hECA3A3134A4ADC25DDDD251D2525DDDC252593936EFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h018A63920092641263F55B1AD24A92491BD392494A92DB64F6F5F5F5F5F5F5F5),
    .INIT_12(256'hFEFEFEFEAD2525934A92DC25DC9349924A4949014A8AD3DC934A4A4A9393934A),
    .INIT_13(256'hFEFEFEFEFEFEF5AC64ADFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEF5F5FEFEFEF6),
    .INIT_14(256'h64ACACABF5FEFEFEFEFEFEFEFEFEFEFFFEFEFD63ACABB4FEFFFFFEFEFEFEFEFE),
    .INIT_15(256'hFEFEF6F6F6F5F5F5F5F66D9249DB92491B6C23DBDB4992D29292DA92242391DA),
    .INIT_16(256'hAE1C65D365AED442929292494949914912ADB5DAACAC23B6FEFEFEFEFEFEFEFE),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hECA3A3894A4A251DDCDD251D2525DDDC1D25DC9325FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h00D36D89001BAC1AACF65B1B924A4A8A1CDBDBDB4A93DBADF6F5F5F5F5F5F5F5),
    .INIT_1A(256'hF5FEFEFEB5651D934A931D25DC934A4A494949014A93D4934A4A014A93938A4A),
    .INIT_1B(256'hFEFEFEFEFDFDF5AC6CFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEF5F5FEFEFEFD),
    .INIT_1C(256'hADACA3F4FEFEFEFEFEFEFEFEFEFEFFFFFFFEB463ACECF4B4F5FEFEFDFEFEFEFE),
    .INIT_1D(256'hFEFEFEFEFEFEFEFEFEFEF69189DB9289236C2392DB5192DAD291DB92242492DB),
    .INIT_1E(256'hFF1C651C1CAE658B8AD3DB92494991491AACF5AC636391ADF5F6FEFEFEFEFEFE),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_043008_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n76 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i42_008,inst_doa_i42_007,inst_doa_i42_006,inst_doa_i42_005,inst_doa_i42_004,inst_doa_i42_003,inst_doa_i42_002,inst_doa_i42_001,inst_doa_i42_000}));
  // address_offset=44032;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFF60073FFFFE0C00DFFFFFFFFFFFFFFFFFC30000067F1B3FFE33C47FF),
    .INITP_01(256'hFFFFFFFFFF007FFFFFE0C00DFFFFFFFFFFFFFFFFFC10000060E1B3FFC23C67FF),
    .INITP_02(256'hFFFFFFFFFB007FFFFFE0C00FFFFFFCFFFFFFFFFFFC1000014001B3FFC62C67FF),
    .INITP_03(256'hFFFFFFFFFF803FFFFFE1800FFFFFFC0FFFFFFFFFFC100001E003B3FF84EC33FF),
    .INIT_00(256'hE3A31B494A93251DDCDD261D2525DDDCDD25DD93DBB7FFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h00246D408964641AF5F55B1B924A001B25D21B244A4A1BF5F5F5F5F5F5F5F5F5),
    .INIT_02(256'hF5FDFEFEB56DDC934A931D25DC934A8A494949418A93934A524A094A9393494A),
    .INIT_03(256'hB5F5FEFEFEFDF5B4ACFEFEF5ACB5FEFEFEFEFEFEFEFEFEFEFEFEACFDFEFEFEFE),
    .INIT_04(256'hAC63ACFEFEFEFEFEFEFFFEFEFEFEFFFFFFFEA2ABECECF4F4F4B5B5B4B4B5F5F5),
    .INIT_05(256'hFEFEFEFEFEFEFEFEFEFFF69291DB9291246CDB92DB9292DBDB91DB9223249224),
    .INIT_06(256'hFFAE1C65D3656EDC93D3DB9249494992D2ACF5AC0088ACF563F5FFFEFEFEFEFE),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hE3A492494ADC25DCDCE5661D2525DCDCDC252594936DFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h001B6D0040D2D2D264645BDB4A4A49631D92236D014964F6F5F6F5F5F5F5F5F5),
    .INIT_0A(256'hF5F5FEFEB56DDC934A93DD25DC8A4A934149414993938B4A4A49498A934A418A),
    .INIT_0B(256'hB5F5FEFEFEFEFDF5ACFEF5ACB5B6FEFEFFFEFEFEFEFEFEFEFEFDB4F5FEFEFEFE),
    .INIT_0C(256'h63ABFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEF4A3ABECECABB4FDFEFEF5F5F5F5F5),
    .INIT_0D(256'hFEFEFEFEFEFEFEFFFFFFFE9291DB91926C24DB92DB9292DBDB49DBDA1B24DB64),
    .INIT_0E(256'hFFFF1C651C1C6E6593D3DB9289494992D263F5ECA4F6FEF5F5F6FEFEFEFEFEFE),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hE41B494A4B252593DCDC66DD2525DCDDDC1D25DC931CFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hD21B920000000000000089924A01D2A41C8964AD0041ADFEF5F6F6F5F5F5F5EC),
    .INIT_12(256'hF5F5FEFEB66DDC8B4A93DD25DC4A4A8A0149499293934A4A4A09494A4A49921B),
    .INIT_13(256'hFEFEFEFEFEFEFEFEACFDF5ADFFF6FEFEFFFEFEFEFEFEFEFEFEBDF5F5FEFEFEFE),
    .INIT_14(256'h63FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFD63ACA3EBAB48DA646C6CBDFEFEFEFE),
    .INIT_15(256'hFEFEFEFEFEFEFFFFFFFFFE9292DB89DA6D1BDA91DA9192DBDB49DBDA23646464),
    .INIT_16(256'hFFFF6E2565DC656EDCD3DBD292494989DA1AECF5F5F6FEFEFEFEFEFEFEFEFEFE),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hA4D28A4A9426DCDB1C1C66DC2525DCDDDCDC25259393B6FFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hACAC1B0000000000000000004A005CA31C896CAD0092B6FEF6F6F6F6F6F6F5EC),
    .INIT_1A(256'hF5F5FEFEB66DDC4B4A93DD25DC4A8A4A41494ADB924A4A4A4909494A4A8A9264),
    .INIT_1B(256'hFEFEFEFEFEFFFEFEF5F5FEB5B6F6FEFEFEFEFEFEFEFEFEFEFEFDF5F5FEFEFEFE),
    .INIT_1C(256'hF4FEFFFFFEFEFEFFFEFEFEFEFEFEFEFEECACACA2EB6B00010000489A6BABABFD),
    .INIT_1D(256'hFEFEFEFEFEFEFEFFFFFFFE9A92DB892364DA9249DA4992DBDB49DBDA236C6C23),
    .INIT_1E(256'hFFFFF71C6E1C65652592DBDA92498949DBD2A4F5F5F5FEFEFEFEFEFEFEFEFEFE),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_044032_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n76 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i43_008,inst_doa_i43_007,inst_doa_i43_006,inst_doa_i43_005,inst_doa_i43_004,inst_doa_i43_003,inst_doa_i43_002,inst_doa_i43_001,inst_doa_i43_000}));
  // address_offset=45056;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFF807FFFFFE1800FFFFFFC61FFFFFFFFFC300001E00133FF8C6C33FF),
    .INITP_01(256'hFFFFFFFFF5C05FFFFFE1010FFFFFFC63FFFFFFFFFC300001E001B7FF096D33FF),
    .INITP_02(256'hFFFFFFFFFEB00FFFFFF3011FFFFFFBC3FFFFFFFFFC302801E006B7FF196919FF),
    .INITP_03(256'hFFFFFFFFFAD007FFFFF2011FFFFFF3DBFFFFFFFFFC303001E006B7FE106919FF),
    .INIT_00(256'h1C924A4A25258BDCDC1C66DC2525DCDDDCDC2525DC8B6DFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hF5F5240000000000000101004A00DB64DC4AADB500DBF6FEFEF5FDF5FEF6ECE3),
    .INIT_02(256'hFDF5F5FEF66E9C4A4AD31D25944A934A410192DB404992934A01494A4A92D264),
    .INIT_03(256'hFDFEFEFEFFFFFEFEFEB5FEFDB4FEFEFEFFFFFEFEFEFEFEFEFEB5FEFEFEFEFEFE),
    .INIT_04(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFDA3ECEC62AB6C0A029B221A9C151412B4),
    .INIT_05(256'hFEFEFEFFFEFEFFFFFFFFAD89D2DA922423929249924992DBDB49DADB24B563AC),
    .INIT_06(256'hFFFFFF6525651C6565DBDBDA92499249D21B12ECF5F5F6FEFEFEF5F5F6FEFEFE),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hDB8A4A9365DC931DDC2525DC2525DC1DDCDC2525DD4B24FFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hF5F51B0000000000414149490092401B1C49B6B50024FEFEF5FEFEFEF5F5ECA3),
    .INIT_0A(256'hFEF5F5FEF66E9B4A4AD32525934A934A4141DB92D2DB929301414A4A4A93D364),
    .INIT_0B(256'hFDFEFEFEFEFEFEFEF5ACFDFEFEFEFEFEFEFEFEFEFEFEFEFEFDACF5FEFEFEFEFE),
    .INIT_0C(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEACACF4ACA2AB1A8900DBB5ADDC145C24F4),
    .INIT_0D(256'hFEFEFEFEFEFEFEFEFFF663D2D292DB64DB9192919249921BDB49D2DB6D6C64FE),
    .INIT_0E(256'hFFFFFFF7DC66DC65651CDBDBD2495149D223915BECF5F5F5FEFEFEF6FEFEFEFE),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h934A4125254A9425932525DC25DDDC1DDCDCDC25259393B7FFFFFFFFFFFFFFFF),
    .INIT_11(256'hF5F62300418A4901494900000024ADD12449F6B5006DFEFEFEFEFEFEF5ECA41B),
    .INIT_12(256'hFEF5F4FEFE6DDB4A8AD42525934A934A01491CD224DB938B01494A4A93D3D364),
    .INIT_13(256'hF5FEFEFEFEF5F5F4ACA3F4FDFDFEFEFEFEFEFEFEFEFDFDFDF5ECECF5FEFEFEFE),
    .INIT_14(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFDACEDF4AB6B64406363236CDBD3939BB5FD),
    .INIT_15(256'hFEFEFEFEFEFEFFFFF563A323919A2323924992499249921BDB4992646C64FEFE),
    .INIT_16(256'hFFFFFFFF256565DC6EDB1B1BD249925192DBDA001BECF5F5F5FEFEFEFEFEFEFE),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h4A01DC259342DCDCDB2525DC25DCDC25DCDCDC2525DC4A6EFFFFFFFFFFFFFFFF),
    .INIT_19(256'hF5FE240093D341490189DB920065F6DA2492F6B600ADFEF6FEFEFEFEECED6489),
    .INIT_1A(256'hFEF5B4F5FE6DDB4A93DC25254B4A9349098A1B64DB4ADC4A014A4A8A93D3DB64),
    .INIT_1B(256'hF5FDF5F5F5ECACABAB63ACF4B4F5F5F5FDFDFEFDF5F5F5F5ACECF4F4FEFEFEFE),
    .INIT_1C(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEF4ACACEBA263DC00ACF56C24DAAD249BB5F4),
    .INIT_1D(256'hFEFEFEFEFEFFFFED5BA3F52348DB24DB494992499289DA239249DBAD63F6FEFE),
    .INIT_1E(256'hFFFFFFFFB6DC6ED36524DB1BDB49929192DBDA49481AA4EDF5F5FDFEFEFEFEFE),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_045056_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n84 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i44_008,inst_doa_i44_007,inst_doa_i44_006,inst_doa_i44_005,inst_doa_i44_004,inst_doa_i44_003,inst_doa_i44_002,inst_doa_i44_001,inst_doa_i44_000}));
  // address_offset=46080;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFF5001FFFFF2023FFFFFF3F3FFFFFFFFFC303001E437B7FE22691DFF),
    .INITP_01(256'hFFFFFFFFFD68013FFFE4027FFFFFF0D3FFFFFFFFFC203001CC77B7FC00C80CFF),
    .INITP_02(256'hFFFFFFFFFDB8010FFFC4007FFFFFFBC7FFFFFFFFFC203409FC7FFFFC04C00EFF),
    .INITP_03(256'hFFFFFFFFFE980003CE0000FFFFFFFFEFFFFFFFFFFE203409CF9FFFF808C00EFF),
    .INIT_00(256'h009225DC01932593DC251CDC25DCDC24DCDCDC25251D9225FFFFFFFFFFFFFFFF),
    .INIT_01(256'hF5FE2400D41C008A0000F66D00ADFEAC6D92F6F600ADFFFEF6FEFDF5F5AD1BD2),
    .INIT_02(256'hFEFEF4F5FE6DDB4A93DC25254A9393490A925B64D393DC01414A4A8ADCD4DC24),
    .INIT_03(256'hF5F5F4ACACECABEBABA3ECF4ECECF4F4F4F4F4F4F5F4F5F4A3ABF4F4F5FEFEFE),
    .INIT_04(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEF5ACECABABA263934A23236C2424F6DBDBB5F3),
    .INIT_05(256'hFEFEFEFEFEFEAC5BA3ECF52300E424924092924992911BDB919124ACB5FEFEFE),
    .INIT_06(256'hFFFFFFFFFF1C6525DC6DDB23DB49929291DB9A499292D21BA4F5F5FEFEFEFEFE),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h93DC934A02DDDC932525DCDC1DDCDCDCDCDC93DC2525DCDBFFFFFFFFFFFFFFFF),
    .INIT_09(256'hEDFEDB8AF71C0092001CFFFFDBADFEFDADDAFEF691B5FEFEFEFEF5F5AC1BDB00),
    .INIT_0A(256'hFEFEF5F5FEB5DB4A93DC25DC429393490989AC6341DDDC00494A4A8BDCD3DC24),
    .INIT_0B(256'hF4ECACECECECECECA3ABF4ECF4F4F4ECECECF4F4F4F5F5ECA3ABACF4ACF5FEFE),
    .INIT_0C(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEACABABA3A2A263D34A92D2641BDB1C00DAB4EB),
    .INIT_0D(256'hF6FEFEFEF4A3A3A4EDF6F6D24924DB4149929289D2DA2392492364B5FEFEFEFE),
    .INIT_0E(256'hFFFFFFFFFFAEDCAED36524DB1B49929292DBD249929ADB1B48D263F5FEFEFEFE),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hDB93490193254ADC1C25DCDCDC93DCDCDCDC93DC25252492B6FFFFFFFFFFFFFF),
    .INIT_11(256'hF5FE246EF765000093AE6D6DB6B5FEFEB61BFEF61BB5FFFEFEF6F6AC1A5B494A),
    .INIT_12(256'hFEFEF5B4FEB5DC4A93DC25DC4A944A490189AC630025DC00494A8A931DD3DC24),
    .INIT_13(256'hECECACECECECECECA3ACF4ECECECECECECECF4F4F4F5F4ACECA3ABECF4ACF5FE),
    .INIT_14(256'hFEFEFEFEFEFEFEFEFEFEFEFEF5A3A3A3A362A2635BD21B5B1A1B92000063F4AB),
    .INIT_15(256'hFEFEF563A3ECECEDAD65DB499224920049924991DBDBDB49DB64ADFEFEFEFEFE),
    .INIT_16(256'hFFFFFFFFFFFFDB6525D3241B2349D2DA92DBD2499292DB239249009264F6FEFE),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h9292494A1D9393DC252593DCDC93DCDCDCDC93DC1D2524926EFFFFFFFFFFFFFF),
    .INIT_19(256'hF5F6DB921CAE6565B6DB00F6FEF5FEFEF623FEF664F6FEFEFEF66C1B64924193),
    .INIT_1A(256'hFEFEFEACFDB51C4B93DD25D34ADC4A490A40AC638A2694004A4A93932594DC24),
    .INIT_1B(256'hECACACECECACECAC63F4F4ECECECECECECECECF4F4F4ABABF4ABABABF4F5ACFE),
    .INIT_1C(256'hFEFEFEFEFEFEFEFEFEFEFEFDAC63A3A262A3A3A2A2A35A5A5A1A1BD11BACACAC),
    .INIT_1D(256'h6C1B00D2ACA45BDB9394DC9292D249494992DB92DBDB929224ACFEFEFEFEFEFE),
    .INIT_1E(256'hFFFFFFFFFFFF6DDBAED3DB1C2449D2DB92DB9249D292DBE39292490048D264AD),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_046080_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n84 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i45_008,inst_doa_i45_007,inst_doa_i45_006,inst_doa_i45_005,inst_doa_i45_004,inst_doa_i45_003,inst_doa_i45_002,inst_doa_i45_001,inst_doa_i45_000}));
  // address_offset=47104;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFED80100000021FFFFFFFFFFFFFFFFFFFE603409C7BFFFF000C206FF),
    .INITP_01(256'hFFFFFFFFFF48030000002FFFFFFFFFFFFFFFFFFFFE600409F07FFFE30082077F),
    .INITP_02(256'hFFFFFFFFFF68030000402FFFFFFFFFFFFFFFFFFFFE600C09FF7FFFC60182037F),
    .INITP_03(256'hFFFFFFFFFFA80300C0006FFFFFFFFFFFFFFFFFFFFE600C09FFFFFF800102037F),
    .INIT_00(256'hDB924ADB9342DCD325259393DC4A25DCD4DC8ADCDC2565DB24FFFFFFFFFFFFFF),
    .INIT_01(256'hF5AC0000001B656DAE006DFFFEFEFEFEFE6CFEFEADF6FEFEF563646C89008AD2),
    .INIT_02(256'hFEFEFEB5F5F6248B9325659393DC4A494A401B1BD32693014A4A939325DCDC25),
    .INIT_03(256'hECACECACECECECA3ABF4ACACECECECECEBECECF4F4ACABA3ABF4ABABACF5F5B4),
    .INIT_04(256'hFEFEF5FEFEFEFEFEFEFEFEF563A3A262A3A3A3A362A2A2591962A3ABACABACAC),
    .INIT_05(256'h00000193938A4B94DDE5DC92924949494A9224DBDBDB51236CFEFEFEFEFEFEFE),
    .INIT_06(256'hFFFFFFFFFFFFFFD366258A1C2491DBDB91DB9249DB92DB2391928A4989490000),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h920093930193D4DC65938B93DC4A25DBDCDC4ADCDC1D2524DBFFFFFFFFFFFFFF),
    .INIT_09(256'hACF5AD64D2000000D324FEFEFEFEFEFEFEADFEFEB5FEFEB56CB5AC4892DB1C64),
    .INIT_0A(256'hB5FEFEFDF5F624939325658ADC93014A4A498A89DC269301524A93932594DC24),
    .INIT_0B(256'hACACACACACABEB63ACB4ABACECACACACEBECECF4ACABECABA3ECF4ABABF4F5F5),
    .INIT_0C(256'hFEFEF5FEFEFEFEFEFEFEF5AB62A26262A3A2A2A3A262A2ABABABABABABACACAB),
    .INIT_0D(256'h49490A4B4B54949DDDE5DC929291494992921CDB24B6246CF6FEFEFEFEFEFEFE),
    .INIT_0E(256'hFFFFFFFFFFFFFF65DC6E8ADB2492DBDB92DA9292DB9223239192924949494949),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h00D38A018A939325254A9393934A2593D4DC4ADBDCDC256D4AF7FFFFFFFFFFFF),
    .INIT_11(256'hACFEFEFEFEB6AD1B496CFEFEFEFEFEFEFEF5F6FEF6FEFEF6FE640000D26565D2),
    .INIT_12(256'hF5F5FEFEF5FE65939325254ADC93494A4A498A8A2525934A524A93D36594DC24),
    .INIT_13(256'hABABABABABEBABA3ECACABEBABABACACABECECAB63ABABEBABA3F4F4ABACF4FD),
    .INIT_14(256'hFEFDF5FEFEFEFEFEFEFDF4636262A3A262A2A2A2A3A362A3A3A3ABABABABABAB),
    .INIT_15(256'h4ADB534A4B949D9DE525DC92D249494A929224DB24FFB5B5FEFEFEFEFEFEFEFE),
    .INIT_16(256'hFFFFFFFFFFFFFFFF8A661D8A24DADBDBDB928992DA9223239192928A49494900),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hD392414A934AD425938A939393922593D4DC4A93DCDC25B64AB6FFFFFFFFFFFF),
    .INIT_19(256'hACF6F6FEFEFEFFFFFEB6FEFEFEFEFEFEFEFEF6FEFEFEFEFEB600000000D29200),
    .INIT_1A(256'hFDF5FEFEF5FE6DDB93252593DC4A4A4A4A4949922525934A524A93DC6EDBDB25),
    .INIT_1B(256'hABABABABABEBA2A3ACACABEBABABACABECECAC6363ABABEBECABABF5F4ABACF5),
    .INIT_1C(256'hFEF5F5FEFEFEFEFEFEF5AB62A3A2A3A36262A2A3A2A3A362A3ABEBABABABABAB),
    .INIT_1D(256'h2525934A93939CDDDDDD9BD3D292499292246DDB6DFEF6FEFEFEFEFEFEFEFEFE),
    .INIT_1E(256'hFFFFFFFFFFFFFFFF25DC6E8A1CDBD3DB92DB8989DB9224234992DA9249494092),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_047104_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n84 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i46_008,inst_doa_i46_007,inst_doa_i46_006,inst_doa_i46_005,inst_doa_i46_004,inst_doa_i46_003,inst_doa_i46_002,inst_doa_i46_001,inst_doa_i46_000}));
  // address_offset=48128;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFB1030180007FFFFFFFFFFFFFFFFFFFFE600C09FFFFFF810202017F),
    .INITP_01(256'hFFFFFFFFFFB1430300007FFFFFFFFFFFFFFFFFFFFF400C09FFFFFF00000201FF),
    .INITP_02(256'hFFFFFFFFFFDB230F0000FFFFFFFFFFFFFFFFDFFFFF000809FFFFFF04000001BF),
    .INITP_03(256'hFFFFFFFFFFD9831F0000FFFFFFFFFFFFFFFF9FFFFF00080FFFFFFE3C000401BF),
    .INIT_00(256'hDB014A924A9325DC41934A934A93254AD4DC4A93DCDCDCB7936DFFFFFFFFFFFF),
    .INIT_01(256'hACF6F6FEF6FEFEFEFFFFFFFEFEFEFEFEFEFEFEFEFEFEFEFE640049484900401C),
    .INIT_02(256'hF5FEF5FEFEF5ADDBDC251CDCDC014A4A4A4900922525934A524ADCDC6DDBD325),
    .INIT_03(256'hABABABABACABA2ABAC63ACABABEBABABACACF56463A3EBABACECABACFDF5ACAC),
    .INIT_04(256'hFEF5F5FEFEFEFEFEF5AC63ECA3A2A3A3A2A262A3A3A2A3A3A3A3ABABABABABAB),
    .INIT_05(256'h25934A4A4B4B5394949493DB9292899292B6B624B5B6FEFEFEFEFEFEFEFEFEFE),
    .INIT_06(256'hFFFFFFFFFFFFFFFFB74A661C8ADBD31C92DBD289DAD224234992DBDBDA899265),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h49498A4A4ADCDC4A928A4A9301DC254A94DC4A4ADCDCDCB72424FFFFFFFFFFFF),
    .INIT_09(256'hACF5F5F5F5FEFEFEFEFFFFFFFEFEFEFEFEFEFEFEFEFEFEF601004000000092D2),
    .INIT_0A(256'hACF5FDFDFEF6AD1CDC25D393934A4A4A4A4A00D3251D93924A4ADCDC6DDBD324),
    .INIT_0B(256'hABABABABACA3A2AB6464A4ABABABABAB64ADADAC63A2ABACACECECABF5FEF5AC),
    .INIT_0C(256'hFEB4F5FDFEFEFEFDF563F5EC62A3A3ABA2ABA3A3ABA2A2A3A3A3ABABABABABAB),
    .INIT_0D(256'h01014B4B0A4A4B4B539393DB92919292DBFFF66DB5FEFEFEFEFEFEFEFEFEFEFE),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFDC1C668AD3D31CDB1BDB91DBD2241B9192DADBDADB256E),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h4A4A4A4AD4DC4A4A9249929201DCDC4A94DC9249DCDC93B76DDBFFFFFFFFFFFF),
    .INIT_11(256'hACF5F5F5F6F6F5FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFF244A49004949248A00),
    .INIT_12(256'hACF4FDFDFEFEAD24924A4A094A4A4A4A4A4A00D325DD93924A92DCDC66DCDB24),
    .INIT_13(256'hABABABABAB62A2AB64AD63A3ABABACAB6C6DDB6DACA3ABECACECF4F4ACFDFEF4),
    .INIT_14(256'hFDB4F5FDFEFEFDF5ACF5F55AA3A2A2ABABA3AB63A2ABA3A3ABABA3ABABABABAB),
    .INIT_15(256'h4A534B535353949C9CDC9BDB9291D2926DFFF66DFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFAE41661C002465DBDB2492DADA241B49D2929224256E25),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h4A494A93934A4A524A4A924A4A1DDC4A94DC9249D4DC8AB7B693FFFFFFFFFFFF),
    .INIT_19(256'h64F5F6F6F6F6F6F6FEFEFEFEFEFEFEFEFEFEFEF5F6FEB6DB92006D6D2424004A),
    .INIT_1A(256'hF4ACF5FEFEFEB52493004A4A4A4A4A49924A49DB25DC93924993DCDC651C1C1C),
    .INIT_1B(256'hACA3A3A3A362A2AB646463A3ABECAB62B6DC926DADABA3ECECECF4F4F4F4FEFE),
    .INIT_1C(256'hF5ACF5FDFEFEF5ACACFEAB63A3A2A2ABECABABAB62A3EBA3A3ABA3A3ABABABAB),
    .INIT_1D(256'h4A934A4B939394949C93DBDA9191DB92B6FFB6F6FEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFD31D6500DB6E24DBD392D2DB241B8992DB6D6E6E6E1C),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_048128_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n84 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i47_008,inst_doa_i47_007,inst_doa_i47_006,inst_doa_i47_005,inst_doa_i47_004,inst_doa_i47_003,inst_doa_i47_002,inst_doa_i47_001,inst_doa_i47_000}));
  // address_offset=49152;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFEDC23E0000FFFFFFFFFFFFFFFF9FFFFF00080FFFFFFFF0000401BF),
    .INITP_01(256'hFFFFFFFFFFECC67E0001FFFFFFFFFFFFFFFFEFFFFF00080EFFFFFDC0000401BF),
    .INITP_02(256'hFFFFFFFFFFF4C67C0181FFFFFFFFFFFFFFFFEFFFFF80080EFFFFFE30000001BF),
    .INITP_03(256'hFFFFFFFFFFF6667C0007FFFFFFFFFFFFFFFFC7FFFFC0081EFFFFFF70006001BF),
    .INIT_00(256'h014A9392494A4A8A494A924A4A25934A93DC8B4A93DC4AB7B792FFFFFFFFFFFF),
    .INIT_01(256'h64F6F6F6FEFEFEFEFEFEFEFEFEFEFEFEF6F6F6F5F5FEADAE1D1CB6B6DB00414A),
    .INIT_02(256'hFEB4ACF5FEF5B56DD301934A4A924A49924989D325DC93924193DDDC65241C1B),
    .INIT_03(256'hA3A3A2A36262A3A3A262ABABABAB62A2ADDC9C25ADACABABECF4F5F5F5F4F5FE),
    .INIT_04(256'hF5ACF5F5FEF5F4ABFEF562A3A2A2A3ABECACA3ECAB62A3EBA3A3A3ABABA3A3A3),
    .INIT_05(256'h4B94530A539394949493DBD29192DBDBFFFFB5FEFEFEFEFEFEFEFEFEFEFDFDFE),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFF6E42651C0025AE24DB92D2DB64DB49DB6EB76E6E6E8A),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h4A4A4A494A4A4A4A0093934A93254A4A93DC8A4A93DC4AB7FF92FFFFFFFFFFFF),
    .INIT_09(256'h64F6F6F6FEFEFEFEFEFEFEFEFEFEFEFEFEF6F5F5F5AC891BAE1C499200898A01),
    .INIT_0A(256'hFEFEACACF5FEF66DDC01924A93934949938A8AD325DC939201DCDCDC252464DB),
    .INIT_0B(256'hABABA3AB62A3ABABACECECABA3A362A3AD241CDC64ADECABABF4F5F5F5F5F5FD),
    .INIT_0C(256'hB4ACF5F5F5F5ACF5FE63A3A3A3A3A3ABECECABABF4AC63A3ECABA3A3ABABABAB),
    .INIT_0D(256'h4B949C0B0A535394DDDCDB9191DB926DFFB5FEFEFEFEFEFEFEFEFEFEFEF5FDFE),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFF8B1C654AD3AE65DB92921B24DB4024B66E6EB72501),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h4949494A4A4A4A4A00DCDC0193DC49929393934A8A934AB7FF93B6FFFFFFFFFF),
    .INIT_11(256'h64F5F6F6FEFEFEFEFEFEFEFEFEFEFEFEFEFEF5F5F5631B00DBD3646DDB494A01),
    .INIT_12(256'hFEFEFEB4ACFDFEB52492924A93934A4A4A8AD2D325D4939201DCDCDC246464D2),
    .INIT_13(256'hABECECECABABECECACAB625AA3AB62ACF66D1C931C6CACF4EBF4F4F5F5F5FDF5),
    .INIT_14(256'hACACF4F5F4ACACFEAC63ABA3A3A3A2A3ECECABA3ECF4ECA362ABABA2A2A3ABAB),
    .INIT_15(256'h94539CDD9CDDE52525E4DB8992DBDBB6F6FEFEFEFEFEFEFEFEFEFEFEFEF5FDFE),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFF658A65DB491DAEDB92922464DA4924B6B6AEB7DC0A),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h8A414A4A494A8A00926E2501DCDC414A9393934A4A934AF7FFDBB6FFFFFFFFFF),
    .INIT_19(256'h64F5F5F6FEFEFEFEFEFEFEFEFEFEFEFEFEFEF5F6F5F5FE6C00B5FFF60092924A),
    .INIT_1A(256'hFEFEFEFEACB5FEFEB524DB4A9393934A4A92DBD31C93934A01E5DC1D1C656492),
    .INIT_1B(256'hA3A3ABABABA2A3A3625AA2EBABA3ACFDF66DDC4ADB6463ECECF4F4F5F5FDFDFD),
    .INIT_1C(256'hABABF4F4ECACF6F663A3A3A3A3A3A3A3ACF4ECA3ABECF5F4AB62A3A3A2A262A2),
    .INIT_1D(256'h9C9C9CDDE5E5DDE5DCDBDB92DA1B6DB5FEFEFEFEFEFEFEFEFEFEFEFEFDF5FDF5),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFF7411D1C89936524919A242492512DB6AEB6B79354),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_049152_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n92 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i48_008,inst_doa_i48_007,inst_doa_i48_006,inst_doa_i48_005,inst_doa_i48_004,inst_doa_i48_003,inst_doa_i48_002,inst_doa_i48_001,inst_doa_i48_000}));
  // address_offset=50176;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFA067C0007FFFFFFFFFFFFFFFFC7FFFFE0285EFFFFFFF0006001FF),
    .INITP_01(256'hFFFFFFFFFFFB067C004FFFFFFFFFFFFFFFFFC7FFFFE0205EFFFFFFE0006001FF),
    .INITP_02(256'hFFFFFFFFFFF9047C099FFFFFFFFFFFFFFFFF87FFFFF0205EFFFFFFE0204011FF),
    .INITP_03(256'hFFFFFFFFFFFDCCFC03BFFFFFFFFFFFFFFFFF8FFFFFF0305EFFFFFFE020E013FF),
    .INIT_00(256'hDC934A414A4A4A00DC6E1C42DC934A8A939393934A9292FFFF24B6FFFFFFFFFF),
    .INIT_01(256'h64F5F5F5FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE6DFEFF1B00DB9393),
    .INIT_02(256'hFEFEFEFEFEACB5FEFEB524939393934A4A921BD31C93934A4A25DC251CAD648A),
    .INIT_03(256'hA3A2A2A2A26262A3A3A3ECABABACF5FEB665D34A932463A2ECECF4F4F5FDFEFE),
    .INIT_04(256'hA3ABF4F4ACB5FFAC63A3A3ABABABA3A3ACF4F4ABA3ACF5F5F4ACA2A2A3A36262),
    .INIT_05(256'h9D9C9D9C9494534A01DCD292DB6D6CB5FEFEFEFEFEFEFEFEFEFEFEFEF5F5FDF5),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFF1C8B65D38ADCDB92DB242491926DB6AEB7B753DD),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hDC93DC4A4A4A4901DB6E254ADC8A4A4A934A93DC930193FFFF65B6FFFFFFFFFF),
    .INIT_09(256'h64F5F5F5FEFEFEFEFEFEFEFEFEFEFEFEFEFEF6FEFEFEF6FEFEFFFF9200DB9393),
    .INIT_0A(256'hFEFEFEFEFEFEACF5FEFEB5DBD393934A4AD21BD3DC9393499225DC251BAD6489),
    .INIT_0B(256'hA3A3A2A2A262ABABABECECABECF5F5FEB6249201936CA362A3ECECF4F5FDFEFE),
    .INIT_0C(256'h63ABECACACFFF563A3A3ABABECABA3A3ABF4F4ACA3A3ECF5F5F4F4ACA3626262),
    .INIT_0D(256'hDDDD9D9D9C949493E423D2DA6DAD6CFEFEFEFEFEFEFEFEFEFEFEFEFEF5F5FDB4),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFAE011D1C8BDBD392DB6C2391DAAEB76EFF6E01DD),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hDC932593004A4900DCB6DC4ADC494A4A934A9325DB00DCFFFF6DB6FFFFFFFFFF),
    .INIT_11(256'h64F5F6F6FEFEFEFEFEFEFEFEFEFEFEF6F5F6FEFEFEFEFEF6FEFFB6004ADB93D4),
    .INIT_12(256'hFEFEFEFEFEFEFEB4F5FEF624DCD4938A49D264D2DB939300D325DD1C63ED648A),
    .INIT_13(256'h63ABABACACA3ABABF4F5F4ECECACF5FE6DDB4A00DCADACA3A2A3ACF4F5FDFEFE),
    .INIT_14(256'h63ABECACF6FEACA3A3A3A3ABECABA3A3A3ECF5F4ABA3A3ECFDFDF5F5F5ECABAB),
    .INIT_15(256'h94DDE5E525E5DD256DDBDA24B5ACB5FEFEFEFEFEFEFEFEFEFEFEFEF5F5F5FDAC),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFD3D31D8AD3D392DB6CE349DBB6B776FF6E0154),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hDC9325934A4A4A0124F71C4A93414A8A9349DB6DDB0024FFFF6DB6FFFFFFFFFF),
    .INIT_19(256'h64F5F6F5FEFEFEFEFEFEFEFEFEFEFEF5ACF5FEFEFEFEFEFEFEFF2400929B93D4),
    .INIT_1A(256'hFEFEFEFEFEFEFEFEB5FEFE24DCDC93924A925C13DB4A9300DC25DD1C64F5648A),
    .INIT_1B(256'hFDF5F5F4AB63ABB4F5F5ACABABECF5FD6D93014A25656CACABA2A3ACF4F5FEFE),
    .INIT_1C(256'h63ACACF6FFB563ABA3A3ABECECACABA3A3ABF5F5ACA3A3A3ECFDF5F5F5F5FDF5),
    .INIT_1D(256'h949C9DDDE5DD25B76DDB24ADF5ACF5FEFEFEFEFEFEFEFEFEFEFEFEF5F4F4F5AB),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFF6D411C651B92921B6CDB4924B7B7B6FF250A95),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_050176_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n92 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i49_008,inst_doa_i49_007,inst_doa_i49_006,inst_doa_i49_005,inst_doa_i49_004,inst_doa_i49_003,inst_doa_i49_002,inst_doa_i49_001,inst_doa_i49_000}));
  // address_offset=51200;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFCCCF803FFFFFFFFFFFFFFFFFF8BFFFFF000DEFFFFFFC020F013FF),
    .INITP_01(256'hFFFFFFFFFFFFCCF80FFFFFFFFFFFFFFFFFFFD3FFFFF8009EFFFFFFC020F033FF),
    .INITP_02(256'hFFFFFFFFFFFFCCF80FFFFFFFFFFFFFFFFFFFF7FFFFFC00FEFFFFFF8000F033FF),
    .INITP_03(256'hFFFFFFFFFFFFC8781FFFFFFFFFFFFFFFFFFFFDFFFFFC00FEFFFFFF0003F873FF),
    .INIT_00(256'hDC932593930192926DFFFF24414A4A92924ADC6EDB006DFFFF6DB7FFFFFFFFFF),
    .INIT_01(256'h63F5F5F5FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFF4A004ADB93DC),
    .INIT_02(256'hFEFEFEFEFEFEFEFFFEB5FE6DDCDC93934A498AD3DB4A52002525DD1CACECA492),
    .INIT_03(256'hF5F5ECA35AABF5FEF5A3A3A3ACF4F5F56D9200DC25DCAE64ABEBA3A3ACF5FDFE),
    .INIT_04(256'hA3ACADF6F6ABA3ABA3A3ABECACABABA3A363ECFDF5A3A3A3A3ECFDF5F5F5F5F5),
    .INIT_05(256'h9C9D9DDDDDDC76FF65246DFEF5ABFEFEFDFEFEFEFEFEFEFEFDFEFEF5ECF4F463),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF6928AAEAE9291246C92512DF7B7F7FFE44B9D),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hDC931D934A499393AEFFFFB6004A4A924A9224B6DB00B6FFFFB6FFFFFFFFFFFF),
    .INIT_09(256'h63F5F5F5F6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFF65004A4AD393DC),
    .INIT_0A(256'hFEFEFEFEFEFEFEFFFEFDB56D25DC94934A4A00939392924125DDDD1CECECA492),
    .INIT_0B(256'hACA3A3ABACF5FEF463A3A3ABECF4F5AC641B9225DCDD6E6DA3ABEBABA3ECF5FD),
    .INIT_0C(256'h63ADF7FFACA3ABABA3A3A3ABACACECECECECACF5FDF4A3A3A3A3ACFDFDF5ACAC),
    .INIT_0D(256'h9CDDDDE525B6FFFF6DB5FEFEACB4FEFEFDFEFEFFFEFEFEFDFDFEF5F4ABF4F462),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF1B1BADAD9291242492926DFFF7FFBFDC4B95),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hDC93DCD4934ADCDCB6FFFFFFDC008A924A9325FFDB00FFFFFFB6FFFFFFFFFFFF),
    .INIT_11(256'h63F5F5F5F5FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFB64A4A494AD394DD),
    .INIT_12(256'hFEFEFEFEFEFEFEFFFEFEFD6D651D94934A4A4193934A0193661D1C1BA3ECA489),
    .INIT_13(256'hACF4F5FDFDF4AC6363A3A3ABECF4F4ABA36CAD25DC25256D63A3ABECECA3ECF5),
    .INIT_14(256'hACB5AEB5ACA3ABA3A3A3ABF4F4F4F4F4F4F5ACACFEFDACA3A3A3A3ACF5FEF5AC),
    .INIT_15(256'h9CDDDDE5B7B7B6B6B5FEFEFDACF5FEFEFDFEFEFFFEFEFEFDFDFDF5ECABF4EC62),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFB5ACF52391926D2492D21BF7FFFFBFD44B9C),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hDC93DCDC93932425FFFFFFFFB792004A8A246DFF9392FFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h63F5F5F5F5F6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFB6498A4A4A4A93D4DD),
    .INIT_1A(256'hF5FEFEFEFEFEFEFEFEFEFEB66D65DC934A414293934900DC261C1BA3A3A36492),
    .INIT_1B(256'hF5F5FDF5AC6363636363A3ABEBECF4A3ABACAC6D6D25DC1C6CA3ABABECF4ABAC),
    .INIT_1C(256'hF66DADACA3ABA3A3A3ABECF4F4F4F4F5F5F5ABACF5FEF5ACABABABABACF5FDF5),
    .INIT_1D(256'hDDDCE5B7FF6E2424F6FEFDF5ACFEFEFDFEFEFEFFFEFEFEF5F5FDF4ABABF4ABAC),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6B4EC6349926DDB92D2C19CF6FFBF93939D),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_051200_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n92 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i50_008,inst_doa_i50_007,inst_doa_i50_006,inst_doa_i50_005,inst_doa_i50_004,inst_doa_i50_003,inst_doa_i50_002,inst_doa_i50_001,inst_doa_i50_000}));
  // address_offset=52224;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFC9B87FFFFFFFFFFFFFFFFFFFFCFFFFFE01BCFFFFFC0103FE77FF),
    .INITP_01(256'hFFFFFFFFFFFFC8F87FFFFFFFFFFFFFFFFFFFFFFFFFFF019CFFFFF80127FEF7FF),
    .INITP_02(256'hFFFFFFFFFFFF99F0FFFFFFFFFFFFFFFFFFFFFFFFFFFF01087FFFE00107FEF7FF),
    .INITP_03(256'hFFFFFFFFFFFF93F9FFFFFFFFFFFFFFFFFFFFFFFFFFFF83003FFF000107FFFFFF),
    .INIT_00(256'hDC93DCDC4ADC256EFFFFFFFFFFFF2400DB6DB6FF4A24FFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hACF5F5F5F5F6FEFEFEFEFEFEFEFEFEFEFEFEFEFFFFB6DB004A924A4A4AD3D41D),
    .INIT_02(256'hACF5FEFEFEFEFEFFFEFEFEFEF66E24DC4A4A4A924A09002526DC1BA3A3A3D201),
    .INIT_03(256'hF4F4ECA36363ECEC6363A3A3A3EBECA3ECAB62ACAD6DDC936DACABA3A3ECF4AC),
    .INIT_04(256'hFFADACABABA3A3ABABACF4ECACACACACB4ACABACACFDFEF5ECECECECACACF4F4),
    .INIT_05(256'h9425FFFFB66E651BF5FDF5ACF5FEFDF5FEFEFEFEFEFEFDF5F5F5ACABABF463F5),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF6F5ACAB2349DB6DD29124A5C153F6F7935394),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hDC931CD34A1C6DB6FFFFFFFFFFFFFF0024B6B6FF496EFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h64F5F5F5F5FEFEFEFEFEFEFEFEFEFEFEFEFFFFB6240000498A934A4A4A93DC1D),
    .INIT_0A(256'hF5F5F5FDFEFEFEFEFEFEFEFEFEF66D1C4A014A4A4A014A2625949263EC640001),
    .INIT_0B(256'hECECA3A2A363A3F5F5ACABABACECABA3ECAC62ABACAD65256564ACABA3A3ECF5),
    .INIT_0C(256'hFFF6A3A3ABA3ABABABABABABECF4F5F5F5F4ECACECF5FEFEF5F4ECF4F4F4F4F4),
    .INIT_0D(256'h8B65F6B66E6E6D64F5F5F4ACF5FEF5F5FEFEFEFEFEFEF5F5F5F4ABABABF4ACF5),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFEF5F5ABAB2300E4649291D2EEE50053AD93538B),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hDC93DC92D325B6FFFFFFFFFFFFFFFFDA6DB6FFFF92B7FFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h8964F5F5F5F6FEFEFEFEFEFEFEFEFEFEFFAE2400004A4A498A934A4A4A93DC25),
    .INIT_12(256'hF5FDF5F5FEFEFFFEFEFEFEFEF5FEB66D9C014A4A4B01D325DC93939324D30053),
    .INIT_13(256'hAB6362A3A3A363F4F5ECF4F4ABABA3ABF4F4AB63F4EDADAD2464ACACABABABAB),
    .INIT_14(256'hFFF5ABABABA3ABABABABACF4F5F5F5FDFDF5ACECF4F5FDFEFEF6F5F5F4F4F4EC),
    .INIT_15(256'h1CA5A465B76EAEADACF4F4ACFEFEF5F5FEFEFEFEFEFDF5F5F5ACABA3ABABACFE),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFB5F5ECABACDA00242489DA645BEDE513814A9393),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hDCDC9349DC6EFFFFFFFFFFFFFFFFFF6CB6B6FFFF24FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h400064F5F6F6FEFEFEFEFEFEFEFEF56CD300004A4A4A4A4A4A4A4A4A4A9CDC25),
    .INIT_1A(256'hACF5FEFEFEFFFFFEFEFEFEFEFDFDFEB6254A4A4A4B011D259302539C9B924A4A),
    .INIT_1B(256'hF4F4F4F4F4F4ABABABACF4F4F4F4F4F4F4F4F4ECACACAC6C6D6DACACACABABAA),
    .INIT_1C(256'hFFACABABA3A3A3A3ABECF4F4F5F5FDFDFEF5F5F4F4F5FDFEFEFEFEFEFDF5F5F4),
    .INIT_1D(256'hFFF75C5CB76EB7FF63ACF4F4FEFDB5FDFEFEFEFEFEF5F5F5F5ACABAB62ACFEFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFEF5F4ABACACD2496DDB491BF6EE0AA4F61441DCB6),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_052224_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n92 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i51_008,inst_doa_i51_007,inst_doa_i51_006,inst_doa_i51_005,inst_doa_i51_004,inst_doa_i51_003,inst_doa_i51_002,inst_doa_i51_001,inst_doa_i51_000}));
  // address_offset=53248;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFF93D9FFFFFFFFFFFFFFFFFFFFFFFFFFFF82001FFA00010FFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFF93F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFC20007C000033FFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000037FFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFF27FFF7FFFFFFFFFFFFFFFFFFFFFFFFFFC000000000067FFFFFFF),
    .INIT_00(256'hD4934ADB24FFFFFFFFFFFFFFFFFFFFB6FFB6FFB66DFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h4A49001BB5F6FEFEFEFEF6B66DDB1C9301934B4A494A4A494A4A4A4A92DCDC25),
    .INIT_02(256'hABECF5FEFFFEFEFEFEFEFEFEFEFEF5FD6D92494A4A4A25DD0A4B4B0A9CDD930A),
    .INIT_03(256'hFEFDF5F5F4AB63ABACF5F5FEFEFEFEFEFDFDF5F5F5B5B4ECECACB6B5ACEBEBAC),
    .INIT_04(256'hF5A3ACABA3A3A3ABECECF4F4F5FDFEFEFEFEF5F4F4F5FDFEFEFEFEFEFEFEFEFE),
    .INIT_05(256'hEDE50194EE6EFFFFADACB5F5FDF5F4FEFFFFFEFEFEF5F5F5F5ABAB63ACFFFFFE),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFF5F4ACABECAC89926DD291ACF5F6ADCA656500D3A4),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h93DCB6FFB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFB6B6FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h8A494900926DF5F5AD65DB920000DCDC4A4A4A4A49494A494A4A4A4A92DC2525),
    .INIT_0A(256'hABABF4FEFEFEFEFEFEFEFEFEFEFEFDF5B51B4A4A019C25930A4B4B534B4B4B93),
    .INIT_0B(256'hF5F5F5F4F4AB63ECF5F5FEFEFEFEFEFEFEFEFEFEFEFDFDF5F5ADF5F5ACECECAB),
    .INIT_0C(256'hACACABABA3ABABABECECF4F5F5FDFEFEFEFEF5F4F4F5F5FEFEFEFEFEFEFEFEFE),
    .INIT_0D(256'hAD53934AA5B6FFFFFE64F5F5F5ECF5FEFEFEFEFEFDF5F4F5F4ABA3ACFEFFFFFE),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFF5ACABABEC6400E36C92D2F5FEF6ADAD5C9265AEF6),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h4A25FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB6FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h4A49494901008A8A0000004A9349DCDC4A4A4A4A494A924A4A4A4A4A93DC2525),
    .INIT_12(256'hABABACF5FEFEFEFEFEFEFEFEFEFEFEFEB524934A01DCDC024B4B53549C944A93),
    .INIT_13(256'hFEFEF5F5F5ABACACF5FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEF5F4ACB4ACEB),
    .INIT_14(256'hABACABABABABABABECF4F5F5FDFDFEFEFEFEF5F4F4F5F5FEFEFEFEFEFEFEFEFE),
    .INIT_15(256'hFFE54A8B13F7FFFFFFADACFEF5ACF6FEFEFEFEFDFDF5F4F4AC63ACFEFEFEFFB5),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFB4ABABECF4230024244863FEFEFEFEB56C24F6FFEE),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h9324FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h014A49014A4A00004A934A939300DCDC4A924A4A4949934A4A924A4A931D25DC),
    .INIT_1A(256'hABABACACF5FEFEFEFEFEFEFEFEFEFEFEFE6DDC4A93DC4A024B4B53549C9494D3),
    .INIT_1B(256'hFEFEFEFEF5ABF5ACADF5FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFDF5B4ACB4EC),
    .INIT_1C(256'hECABABABABABABACECF5F5F5FDFEFEFEFEFEF5F5F5F5F5FEFEFEFEFEFEFEFEFE),
    .INIT_1D(256'hFFEE41D3C1EEFFFFFFFF6CF5ACB4FEFEFEFEFEFDF5F5F4F4ABACFEFFFEFEFE6C),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFACABABF4ECDB4924DB48ADFEFEFEFEF56CFEFFA509),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_053248_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n100 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i52_008,inst_doa_i52_007,inst_doa_i52_006,inst_doa_i52_005,inst_doa_i52_004,inst_doa_i52_003,inst_doa_i52_002,inst_doa_i52_001,inst_doa_i52_000}));
  // address_offset=54272;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFF27FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000067FFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFF6FFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000067FFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFF4FFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000C7FFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFF4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000C7FFFFFFF),
    .INIT_00(256'h9325B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h414A49014A4A4A4A8A9301529301DCDC4A934A4A4941939301934A4A93252693),
    .INIT_02(256'hECECECACACF5FEFEFEFEFEFEFEFEFEFEFEF66593524B4B534B4B53949C93938A),
    .INIT_03(256'hFEFEFEFEF5F5FEB5FEB5FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFDF4ACAC),
    .INIT_04(256'hECABABABABABABACF4F5F5FDFEFEFEFEFEFEF5F5F5F5F5FEFEFEFEFEFEFEFEFE),
    .INIT_05(256'hB5FF94428B5BF6B7BFFFF6ACACF5FDFEFEFEFEFDF5ECECACACFEFFFFFFFEB4AC),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFEACABECF4AC92922491DAFEFEFEFEF5F5FEFFF6524A),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hDC25B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h4A4A49494A4941494A8A0192930193DC4A924A4A4901939301934A4ADC25254A),
    .INIT_0A(256'hACECECECECF4FDFEFEFEFEFEFEFEF5F5FDFEB6DC4A4B4B9494540B4B934A0901),
    .INIT_0B(256'hFEFEFEFEF5F5FEB5FEB5FEFEFEFEFEFEFEFEFEFEFEFFFFFEFEFEFEFEFDFDF5AC),
    .INIT_0C(256'hABABABABABABACECF5F5FDFEFEFEFEFEFEFEFDF5F5F5F5FEFEFEFEFEFEFEFEFE),
    .INIT_0D(256'h5BFFEE01D34AD26DFFFFFFB563F5FEFEFEFEFEF5F5ECECACF5FFFEFFFFFEABF4),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFEACABF4F4AC491B24006CFEFEFEFDB4FEFEFEF6938B),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hD46D6EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h4A4A49414A4949498A92018AD34193DC938A4A494A498ADB4A924A93256EDC01),
    .INIT_12(256'hECECECF4F4F4F5FEFEFEFEFEFEFEFDF5F5FDFE6DDB53534B94DDDD9C4A094A4A),
    .INIT_13(256'hFEFEFEFEF5ACFEF6ADF5FEFEFEFEFEFEFEFEFEFEFEFFFFFFFEFEFEF563ACACEC),
    .INIT_14(256'hABABABABABABACF4F5F5FDFEFEFEFEFEFEFEFDF5F5F5F5FEFEFEFEFEFEFEFEFE),
    .INIT_15(256'h4AEDFFA40A0ACA64F7FFFFFFB6ADB5F6FEFEFDF5F4ACACACFFFFFEFEFEADACEB),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFE6BACF4F4634924DB00B5FEFEFEF5F5FEB6B6FF9C8A),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h93256DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h4A4A49414A4A494A4A93014AD34A8BDC93934A494A4A4ADC934A4A93256E934A),
    .INIT_1A(256'hABACACF4F5F5F5F5FEFEFEFEFEFEFEFDF4F5FEF625DC9494949CDDDD9CE49301),
    .INIT_1B(256'hFEFEFEFEF5ABFDFEF6F5F5FEFEFEFEFEFEFEFEFEFEFFFFFFFEFEF463A3A363A3),
    .INIT_1C(256'hABABABA3ABABECF4F5F5FDFEFEFEFEFEFEFEFEF5F5F5F5FEFEFEFEFEFEFEFEFE),
    .INIT_1D(256'hD353FFFF5C53F6AD13EEAE76FFFFF7F6B6B5B5AC6C632364FFFFFEFEFDACF4EC),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFF66BECF4AC23492492D2FEFEFEFEF5FDF6F6FEFE9B52),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_054272_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n100 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i53_008,inst_doa_i53_007,inst_doa_i53_006,inst_doa_i53_005,inst_doa_i53_004,inst_doa_i53_003,inst_doa_i53_002,inst_doa_i53_001,inst_doa_i53_000}));
  // address_offset=55296;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000C7FFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFE5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000183FFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFE9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000183FFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFCC000000303FFFFFFF),
    .INIT_00(256'h932525B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h4A4A49494A4A4A4A934B014ADB4B4ADC93934A494A4A4AD3934A4ADC6E254A93),
    .INIT_02(256'hA3ABACF4F5F5F5F5FDFEFEFEFEFEFEFEF5ACF5F5B56D25DD9CDCDC9C9CDD5201),
    .INIT_03(256'hFEFEFEFEF5ABF4FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFEFEB463A3A3A3A3A3),
    .INIT_04(256'hABABABABABECECF4F5FDFEFEFEFEFEFEFEFEFEF5F5FDFDFEFEFEFEFEFEFEFEFE),
    .INIT_05(256'hD309A4F6ADF6F61AA4F66DB6F7FFFFFFFFFFFFFFF6AE6D6DB6FFFFFEACF4F4AC),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFF5ABF4F4AC1A92234024FEFEFEFEF5FEB5F6FEF6A45A),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h93DC25B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h4A4A49494A4A4A4A934A0149DC93099393934A498A4A4A9393934A256E934A93),
    .INIT_0A(256'hABABACF4F5F5FDFDF5FEFEFEFEFEFEFEFEF5ACF5B56C6E26DDDDDC93DDDD4A49),
    .INIT_0B(256'hFEFEFEFEFDACACFDFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEB462ABABA3A3A3A2),
    .INIT_0C(256'hABABA3ABABACF4F5F5FDFEFEFEFEFEFEFEFEFEFDFDFDFEFEFEFEFEFEFEFEFEFE),
    .INIT_0D(256'h8A53121BB5FEEDACFEFE5CAEFFFFFFFFFFFFFFF7B7B6B76EB6FFFFF5ACF4ACAC),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFF5ACF4F4ACD2DB1B40B5FEFEFEFEFDFEB5B6F6F5F59B),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h93D4256EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h4A4A49498A4A4A4A934A4941DB93019393934A494A8A4A8A9393936E240193D4),
    .INIT_12(256'hABABECF4F4F5F5FDFDFEFEFEFEFEFEFEFEF5ACACACADB76E26E5DC9CDDE54A49),
    .INIT_13(256'hFEFEFEFEFDF4A3F5FDFDFEFEFEFEFEFEFEFEFEFEFEFEFEAC63ABABACACABABA3),
    .INIT_14(256'hABABABABABECF4F5FDFEFEFEFEFEFEFEFEFEFEFEF5FEFEFEFEFEFEFEFEFEFEFE),
    .INIT_15(256'hE3ECEDF5F5F5ECF5FEF55B0AEEFFFFFFFFB7B66E6EB66E76FFFFFEACF4F4ECAC),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFB5ACF5F46C911BD2DAF5FEFEFEFEFEFEFEB5F6F6ECA3),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h9393256DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h4A4A4A498A4A4A4A934A490193D40193939392494A934A4ADC93256D4A4A93DC),
    .INIT_1A(256'hABABACF4F4F5F5FDFDFEFEFEFEFEFEFEFFFEF5AB63F6FF6E2626E5E626254949),
    .INIT_1B(256'hFEFEFEFEFEF4A3F4FEF5F5F5FDFEFEFEFEFEFEFEFEFE6C001AA4ABABACACACAB),
    .INIT_1C(256'hABABABABACF4F5F5F5F6F6FEFEFFFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_1D(256'hF4F5F5F5ECACF5F5FEED120153ADFFF7B66DAEAEAE6E76FFFFFFF5ACF4ECECAB),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFACF4F5F56492DB9123FEFEFEFEF6FEFEFEFEFEFEF6ED),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_055296_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n100 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i54_008,inst_doa_i54_007,inst_doa_i54_006,inst_doa_i54_005,inst_doa_i54_004,inst_doa_i54_003,inst_doa_i54_002,inst_doa_i54_001,inst_doa_i54_000}));
  // address_offset=56320;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFE3FFFFFE1FFFFFE0FFFFFFFFFFC3FFFFFFF88000000201FFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFE3FFFFFFE07FFF003FFFFFFFFF81FFFFFFF80000000601FFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFE7FFFFFFE0FFFF001FFFFFFFFF00FFFFFFFC0000000401FFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFC7FFFFFFFCFFFE0007FFFFEFFE007FFFFFFE0000000800FFFFFFF),
    .INIT_00(256'hD493DC25B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h4A4A4A014A4A4A4A934A490193DC4A929393924A4A934A9393936E93008A93DC),
    .INIT_02(256'hAB63ACF4F4F4F5FDFDFEFEFEFEFEFEFEFEFEFDACACFFFF6E25DCDDE626E54A49),
    .INIT_03(256'hFEFEFEFEFEF5ABACFEFDF5F5F5FDFEFEFFFEFEFEFF6C004900D2ABABACB4ECEC),
    .INIT_04(256'hABABABACAC6C23DAD29292DA6CF6FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_05(256'hACF5F4ECACECEDEDF5F65BC9C180CA1B64ADAEAE6D6DFFFFFFFEACF4ECECECAB),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFACF5F5F523D2DB896CFEFEFEFEFEFEFEFEFEFEFEFEF5),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hDC93DC25B6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h4A4A4A014A4A4A4B934A490193DC4A4A93934A4A4A934A934A252500498A93D4),
    .INIT_0A(256'hA363ABF4ECF4F5F5FEFEFEFEFEFEFEFEFEFEFEACFEFFFFB665DC4B549C9C9341),
    .INIT_0B(256'hFEFEFEFEFEF5EC63F5FEF5F5F5F5FDFEFEFEFEFE6C00494A4A00D2ABACACB4F4),
    .INIT_0C(256'hABA3A363D20000000000000000496CFFFFFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_0D(256'hFEECACF5F5EDACEDFEADAC63A4A41340CAD3D3DCD3B6FFFEFFF5ACF4ECECABAB),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFACF5F5B523DA9AD1ACFDFEFEFEFDFEFDFDFDFEFEFEFE),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hDC9494256DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h4A8A4A014A4A4A4B934A494993DC934A93934A4A4193924ADC25934A004A9393),
    .INIT_12(256'hF563A3ECECF4F5F5FEFEFEFEFEFEFEFEFEFEB5B6FFFFFFFF6E25DC5353E5DC01),
    .INIT_13(256'hFEFEFFFEFEFDF41AADFEF5F5F5F5F5F5FEFEFEAD00494A010A5301D2ACECACF5),
    .INIT_14(256'hA262631A00004949494949494900001BFEFFFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_15(256'hFEF6ADF6ECACECF5ED63ADF6FEF61B408181410024FFFFFFFEACECF4F4EBABA3),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFEACF5F4B51BD2911AACF5FEFEF5F5F5F5F5F5F5F5F5F5),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hDCDC93DC25FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h8A8A4A414A4A4A93934A49494ADC934993934A4A4193934A25DCDC9249499393),
    .INIT_1A(256'hF563A3ECABF4F5F5FEFEFEFEFEFEFEFEFEB5B5FFFFFFFFFFF76525DDE5E5944B),
    .INIT_1B(256'hFEFFFFFEFEFDF5D223FEFDF5F5F5F5F5FDFDB500004A4B93534B544ADAACACAC),
    .INIT_1C(256'hA2A21A4040494909010000004149490091B5FEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_1D(256'hF5FEB56CECECECECACEDF6FEB56D655C530A8989F6FFFEFFF5ACF5ECABA26363),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFF6ACF5F5F5DB929122ACF4F5FEF5F4F4F4F4F4F4F5F5F4),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_056320_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n100 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i55_008,inst_doa_i55_007,inst_doa_i55_006,inst_doa_i55_005,inst_doa_i55_004,inst_doa_i55_003,inst_doa_i55_002,inst_doa_i55_001,inst_doa_i55_000}));
  // address_offset=57344;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFC7FFFFFF7FFFFC0003FFFFE7FC003FFFFFFE0000000000FFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFCFFFFEFC01FFF80001FFFFE7FC003FFFFFFF0000000000FFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFEFFFFE7E03FFF00000FFFFE7F8000FFFFFFFA0000000007FFFFFF),
    .INITP_03(256'hFFFFFFFFFFFEFFFFE0FFFFFE000007FFFE3F80007FFFFFFC0000000007FFFFFF),
    .INIT_00(256'h94DC94DC25B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h4A524A014A4A9253934A494A4ADC934993938B4A019393DC9393DD934A494A93),
    .INIT_02(256'h6564ABABA3ACF5F5FDFDFEFEFEFEFEFEF5B5FFFFFFFFFFFFE453ADE5DDDD9453),
    .INIT_03(256'hFFFEFEFEFEFEF5D1D2FEFEFDF5F5F5F5F5FEDB00934A014A939353534BDC6E6D),
    .INIT_04(256'h631B00000909494900004101010149490049B6FFFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_05(256'hF4F5AC23ACF5ACECECF5F55C81135C6465651C6DFFFFFFFEACEBAB63A3A2A2A2),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFF5B5FDF5B5DB52D163ACECF5F5F4F4F4F4F4F4F4F4F4B4),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h94DCDC941D6EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h4A934A014A4A9393934A494A4ADCDC498A938B4A499293939393DD944A4A4993),
    .INIT_0A(256'h6D6CECEBA2ABF4F5F5FDFEFEFEFEF5ADB5FFFFFFFFFFFFED534A656E9C9C944B),
    .INIT_0B(256'hFEFEFEFEFEFEF59100B6FEFDF5F5F5F5FD6C004A5393934B024B9393934A256E),
    .INIT_0C(256'h23490049094A4A010001010101010101490049B6FEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_0D(256'hF4B564D263ACA4F5F5A4D140818180818A8A8AFEFFFEFFF563A262A3A3A2A2A3),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFF5B5FDF5B5DB0919A3ACACF4F4ACF4F4F4F4F4F4F4F4F4),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hDC94DCD4DC25FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h4B8A8A414A4A9393934A494A4ADCDC4A4A938B4A494A93499393DCDC4A4A498A),
    .INIT_12(256'h6EF6B4ACA362ACF4F5F5F5B5B5ADADB6FFFFFFFFFFFFED524A9CF6AE259C2594),
    .INIT_13(256'hFEFEFEFEFEFEF589006DFEFDFDF5F5F4F591004A0A539494944A4A93949493DC),
    .INIT_14(256'h4A0049090A024A01014949090901010100490000B5FEFEFEFEFEFEFEFEFEFEFE),
    .INIT_15(256'hF4F52489D2246464B5B51BD281804040400064FFFEFEFFFE6362A3A2A3A26323),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFF5F5F5F5B51B005AABACACF4F4ACF4F4F4F4F4F4F4F4F4),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h93DCDCD4DC25B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h9C938A494A4A8B93934A4A4A4AD4DC4A4A938B4A4992DC4A9394DCDC8B8A9201),
    .INIT_1A(256'h9325646CAC6363ACACACACB5B5F6FFFFFFFFFFFFFFED524A53F6E552F62EDDE5),
    .INIT_1B(256'hFEFEFEFEFEFEB64900DBFEFEFEF5F5FD2300494A0A0A4B949C9C944B4B949C94),
    .INIT_1C(256'h014A010A024A4A010A0A0A090901090000004900006DFFFEFEFEFEFEFEFEFEFE),
    .INIT_1D(256'hF4B5235192D2D292B5FEF6F5EDADAD64646CFFFFFEFEFEFFFEAB62A2A2A32340),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFF5F5F5F5F51B00A3ACACECF4ECACF4ECF4F4F4F4F4F4EC),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_057344_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n108 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i56_008,inst_doa_i56_007,inst_doa_i56_006,inst_doa_i56_005,inst_doa_i56_004,inst_doa_i56_003,inst_doa_i56_002,inst_doa_i56_001,inst_doa_i56_000}));
  // address_offset=58368;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFEFFFFE0FFFFFC000003FFFE3F00000FFFFEFC0002000203FFFFFF),
    .INITP_01(256'hFFFFFFFFFFFEFFFFE07FFFF8000000FFFE3E000007FFFFFE0002021303FFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFE07FFFF00000001FFE1E000001FFFB7F0002004303FFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFE0FFFFE000000003FE1C000007FFEFFF8000000181FFFFFF),
    .INIT_00(256'h4ADCDCDCD4DCAEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hDD9C52494A4A9393934A4A4A4A931D8B498A924A4992DC9393DC94DD934A1C93),
    .INIT_02(256'hDD9493DC256DADADADB6F7FFFFFFFFFFFFFFFFFFA54A93C1EDEE4A8AA4BF9C94),
    .INIT_03(256'hFEFFFFFEFEFEB5000048B5FEFEFEFEAC00000141494A0A4B9494DD9C534B949D),
    .INIT_04(256'h490101424A4A09010A0A0A4A014141000000004900006CFEFEFEFFFEFEFEFEFE),
    .INIT_05(256'hF4B4239189D292481AF5ACACF5FEFEFEFEFFFFFFFEFEFEFEFFFEAC6263634900),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFADF5F4F5F51B91ABACACF4F4ACACECACF4F4F4F4F4F4EC),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h00D3DCDCDCDC6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h9DE593014A4A9393934A4A4A4A931D94414A8A4A498A1C934ADC931DD4012525),
    .INIT_0A(256'h9DDDDD9C9C256D6EB7B7B7B7B7BFBFBFFFFFEE5C024A4AE5EE53934AEDFFBFDC),
    .INIT_0B(256'hFEFEFEFEFEFF6D0009006CFEFEFEF69200490101494A4A0A4B93935393490193),
    .INIT_0C(256'h00014A4A8B4A010A0A0A4A010149010049090001490100DA6CB5FEFEFFFEFEFE),
    .INIT_0D(256'hF4B4239189929291D1ABACACF5FDFDFEFEFEFEFEFEFEFEFEFEFEFEFE63400049),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFADF4F4F5F51ADAECACECF4F4ACECECABECF4F4F4F4F4EC),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h9300DCDDDCDC24FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h53DDE54A49499393934A4A4A4A921DD4014A8A4A4A8ADC93011C93DDDC0124B7),
    .INIT_12(256'h53949CDD9C02DC6E2E6E6EB6B7B7B6B6E59C0A0A01C1EEF6C1424A9BFFFFFFB6),
    .INIT_13(256'hFEFEFEFEFEFF6D004A00DBFEFEFE23004A4A4901090A0A4A4A4A010000000101),
    .INIT_14(256'h014A9393934A010A0A0A0901494900094A4A4A09019393010000DB6CB6FFFFFF),
    .INIT_15(256'hF4B423929192DA91D1ABABECF5FDF5FEFEFEFEFEFEFEFEFEFFFEFEFE92004900),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFEACF4F4F4F51A23ECECECF4F4ACECEBABECF4F5F4F4F4F4),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h6D00D4DDDCDCDCB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h770A9CDC49498A93934A4A4A924ADDDC014A4A4A4993DCDC00DCDCDCDD4A92B7),
    .INIT_1A(256'h024B9393001C65666E6EAEADADA55C134A530AC113A5EE5C010153EDFFFFFFFF),
    .INIT_1B(256'hFEFFFFFEFFFF6D014A0049B6FF6C004A4A0A4A4A0109094A4A01494900000909),
    .INIT_1C(256'h4B9394934A010A0A0A09014A4A01014A4B4B4B0193939394944B000049DB6DB6),
    .INIT_1D(256'hF4F523D29291DB921AABABF4FDF5F5FEFEFEFEFEFEFEFEFEFFFEB59100490009),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFEACECF4F5F41A64F4ECF4F4F4ACECEBABACF4F5F4F4F4F4),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_058368_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n108 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i57_008,inst_doa_i57_007,inst_doa_i57_006,inst_doa_i57_005,inst_doa_i57_004,inst_doa_i57_003,inst_doa_i57_002,inst_doa_i57_001,inst_doa_i57_000}));
  // address_offset=59392;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFE0FFFFC0000000007C18000007F8FFFFC000000981FFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFE1FFFF0000000000000000200001FFFFE0010029C9FFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFE9FFFF000000000000000030001FFDFFF0010028C8FFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFE9FFFFC000000000008000701FFFFFFDF8010120E4FFFFFF),
    .INIT_00(256'hFF9301DDDDDCDC6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFF764BDC93418A93934A4A4A924ADCDD494A4A4A4993DCDC00DCDCD4259300B7),
    .INIT_02(256'h4A010100926425251C1B1B130AC1C1C152521264655C0A934A0AEDF6FEFFFFFF),
    .INIT_03(256'hDB6CB6F6F6B6DC939301006DB600004B534A4A4A090909494A4A000009090149),
    .INIT_04(256'h9494944B09094901014A4B4A01094A4B54930A53949353549494934900000049),
    .INIT_05(256'hF4F523DAD2499B9263ABECF5F5F5FEFEFEFEFEFEFEFEFEFFFE24000000005353),
    .INIT_06(256'hFFFFFFFFFFFFFFFFF6ACECF4F5F41AACF4F4F4F4ECACECACA3ACF4F5F5F4F4F4),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFF6D01D425DCDC25FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFF6E939C0A4A93934A4A4A934ADC1D4A494A4A4993DCDC00DB259425DC016D),
    .INIT_0A(256'h49014949498A41414140414081C1C154A45BF66D65130193525BF5FEF6FFFFFF),
    .INIT_0B(256'h00000001014A4B9494930152528B934B4B4B4B4A4A494949018A1C8A010A0149),
    .INIT_0C(256'h9494934A010101014A934B014A4A5354944A4A9C930A949494944A00494A0100),
    .INIT_0D(256'hF4F463DADA49921B6CACF5F5F4F5FEFEFEFEFEFEFEFEFFB5490000014A939494),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFF5ACECECF5F462ACF4F4F4ECECACECACACACF4F5F5F5F4AC),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFF934A1DDDDCDCB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hF7FFFF6E9C4A4A93934A4A4A934ADC1D8A414A494993DCDC009325931DDC01DC),
    .INIT_12(256'h010100004992938ACAD2D31C5C65A5F7AD64FF6CADF6C052A3A3F5FEF6F7F7F7),
    .INIT_13(256'h4A494A014A9494539393934A539494534B9393534B41014A00D2A45B00090141),
    .INIT_14(256'h94534A00004A4B9393534A4A4B53949493014A4A01939C4B94930001094A4A49),
    .INIT_15(256'hF4B423D223914863ACF4F4F4F5FEFEFEFEFEFEFEFEFEFFB5DB004A939C949494),
    .INIT_16(256'hFFFFFFFFFFFFFFFFB4ACACACF5AC63F5F4F4F4ECECACACADADACB4F5F5F5F4AC),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hB6FFB6009325DDDC6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h135B64AD1C934A928A8A4A4A938ADC2593014A494A93DC1D018A2593DDDD4B93),
    .INIT_1A(256'h01004964AE656565656565656D656564F5ADFEF5F5F6A3A3ECE3F4F6AD1BCA0A),
    .INIT_1B(256'h014B93534A9CDCD31C49494A4B949C9C934B939494534A090012E39B80000141),
    .INIT_1C(256'h4B010049939494944B0A4A539494949309014A025394944B9201004A934B0101),
    .INIT_1D(256'hACB463D22391D1ACECF4F4F4FDFEFEFEFEFEFDFDFEFEFFFFFF64939D9D959493),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFACABABACF4AC63F5F5F5F4ECECACADADAEADF4F5F5F5F5F4),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_059392_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n108 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i58_008,inst_doa_i58_007,inst_doa_i58_006,inst_doa_i58_005,inst_doa_i58_004,inst_doa_i58_003,inst_doa_i58_002,inst_doa_i58_001,inst_doa_i58_000}));
  // address_offset=60416;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFEBFFFFE00000000001C000707919FFFC68010120E2FFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFEFFFFFE00000000003C00070FC1DFFFFFC010124F27FFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFEFFFFFF60380000003E00078FC0DFFFFFF010124FB7FFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFEFFFFFFF03C0000003F001FFFFFFFFF80F810114797FFFFF),
    .INIT_00(256'hB6FFFFDC01DD25DC24FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hCA130AC112D28A8A934A4A4A9392D32593014A494A93DC1D4A4925DCDCDD9301),
    .INIT_02(256'h4924ADF5F6D3CA0AD3CAD36D1B40811BF6ADFEF6F5FEF4ACF5ECF4F5AD5CCA81),
    .INIT_03(256'h4B9494530193D35CA41B00014A549C9C9C9353939494934A001BA3A3D1004900),
    .INIT_04(256'h000153949494944B4B5393949595944A01014A939494934A00014A94944B0101),
    .INIT_05(256'hABAC63D223D163ECF4F4F4F5FEFEFEFEFEFDFDFEFEFEFEFEF5F625539D948B4A),
    .INIT_06(256'hFFFFFFFFFFFFFFFFACABABACF4AB6BF5F5F5B4ACACACACADADACF4F5F5FDF5EC),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h6DFFFFB741D425DCDCB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hE5E5EEE5E45B418A4A4A4A4A93939325D4014A494A93DC1D4A0124DCDC259401),
    .INIT_0A(256'h24ADA363ED5B80C1C18940ACF65280E4F6F5FEF6F5F5FDACECF5ECF5F6F6EEEE),
    .INIT_0B(256'h9494945301491BA3A3A3D1004A53949C9D94535394949493005BA3A3DA000000),
    .INIT_0C(256'h92939C94945301010A93949CDC944A01024A939C9C944B014A9394944B4A014A),
    .INIT_0D(256'hECAC63DA1A63ACF4F4ECF4FEFEFEFEFEFDFDFEFEFEFEFEFEB4FEFFDC534A0100),
    .INIT_0E(256'hFFFFFFFFFFFFFFFEACABABACF463ABFDF5F5F4ACABECAC6CACACF5F5F5FDF5F5),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h24FFFFFF254A1D25D46EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h9CA4EDF6F7F6EEAEDC01934A93D49325DC414A0192DCDC254A0024DC9325DC01),
    .INIT_12(256'hACA35A62ECA4808180800089F5EC80EDF5F5FEF6ACECF5F5ADF6F6ADADA4A49C),
    .INIT_13(256'h9C9C944B0A001AA3A3A363894A5394D49DDD935394949393D363A3A31B0049DB),
    .INIT_14(256'h939C9494540125B6AEDCD3DC930101014A94949D944B0A939C9494934A014A93),
    .INIT_15(256'hEBAB63DA1AACF5F4ECF4F5FEFEFEFEFEF5FDFEFEFEFEFEFEB4F5FE6D93242DE4),
    .INIT_16(256'hFFFFFFFFFFFFFFF6ACABABACAC63ACFEFDF5F4ECECF4F4ACB5F5F5F5F5F5F5F5),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h93FFFFFFF74BD425DC24FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h8080404013A5F6F7AE8B4A8A93DC4B25DC4A4A0093DCDC254A00DC259325DC4B),
    .INIT_1A(256'hAB6262A2A3ADA5A4A4646464ADF563F5F5ADF6F5A3ABECF5F6FEFFAD6480C0C0),
    .INIT_1B(256'h9C9C9453014963A3A3A3631B4A4B94D4959494935394941CA4A4E3E3631B6D65),
    .INIT_1C(256'hDD934B4B01DCFFFFFFB6DB8A4149094A939C9D94534B949C9494945309095394),
    .INIT_1D(256'hEBA363D163F4F4ECACF4FDFEFEFEFEF5F5FEFEFEFEFEFEFEB4F5FE6D2424242D),
    .INIT_1E(256'hFFFFFFFFFFFFFFF6ECABABACAC62F5FEFDF5ACECACF5F5F5F5F5F5F5F5F5F5F5),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_060416_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n108 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i59_008,inst_doa_i59_007,inst_doa_i59_006,inst_doa_i59_005,inst_doa_i59_004,inst_doa_i59_003,inst_doa_i59_002,inst_doa_i59_001,inst_doa_i59_000}));
  // address_offset=61440;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFF1E7F0000007F0E7FFFFFFFFFBF1C101147DBFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFE0FFF8000387F9FFFFFFFFFFF3FF2101147CBFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFE0B7FF1807FFFFFFFFFFFFFFE3FFC181107EDFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFE0F7BFFC0FF7FFFFFFFFFFFFD3FFE183123E5FFFFF),
    .INIT_00(256'h01B7FFFFFF6D4A1D26D4B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h65241C13C1C1C193DC538A4A93DC4A25DC4A4A0093DCDC254A01DC259325DC94),
    .INIT_02(256'hA362A2A3A2A3ECF4F5F5FEFEECECECECF5ACECF4ECA3ECECF5FEFE6D25DC6EAE),
    .INIT_03(256'h939494530064AD5BA3E3E3A3D2014A8B125B5BCA401BA4ECECECECECACAC6463),
    .INIT_04(256'h2C241CDB006EFFFFFFF6631A0001539C9D9C9C534B9C9D9C9494934A0141D3D3),
    .INIT_05(256'hABA3625AECF4F4ACF4F5FEFEFEFEFDF5FDFEFEFEFEFEFEF5ACF5FE23DB924924),
    .INIT_06(256'hFFFFFFFFFFFFFFF5ECABABACAC63F5FDF5F5ACACACF4F5F5F5F5F5F4F4F4F5F4),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h016EFFFFFFFFDC9426DC65FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hF6F6AEAEEDE5E49CCACA138A93DC4A25DC4A4A00DCDCDC254A01DB259325DC94),
    .INIT_0A(256'h62A3ECF4AC6362A3ABF4F5FEF5ACECECF5ECECECECEDACECF5F5B624D3DCAEF6),
    .INIT_0B(256'h1BD3930ADC6DAD63A4E3E3A363D2921CACECA41B5BEDF5ECF4ECECECECA4635B),
    .INIT_0C(256'h2464656D246EFFFFFFAD63A31BD393D4DC949341D3DC9C9C9494534A0089645B),
    .INIT_0D(256'hABA362ABF4ECACF4F5FDFEFEFEFDF5F5FEFEFEFEFEFEFEF5ACFEFEDADB9292DB),
    .INIT_0E(256'hFFFFFFFFFFFFFEF5ECABABAC6363F5FEFDF5ACABF4F5F5F5F5F5F5F4ECF4F4EC),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h0124FFFFFFFF6E422525DCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h6CA4A464ACA4EDF6F6648A8293DC0125254A4901DCD4DD254A4A932593DDDDD4),
    .INIT_12(256'h62ACF4F5F5F4AB62A3A3ECF5FEACACA3ECECECECF5F5F6F6B56C6DDC93D31BAC),
    .INIT_13(256'hA3A46D252524AEA4A4E3E3E3A4A4A4EDECF4ECECF5F5F5F4F4F4F4F4F5AC631A),
    .INIT_14(256'h23DB2424DB24FFFFFF2464A3A3A41B13D3D2895B64DB949C94934A49001BA3A3),
    .INIT_15(256'hABA3A3ECF4ACACF5FDFEFEFEFEF5F5FDFEFEFEFEFEFEFEB4ACFEFE92DBD292DB),
    .INIT_16(256'hFFFFFFFFFFFFFEF5F4ABABAB6363F6FEFDF5ACABF5F5F5F5F5F5F5F4ACACECEC),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h4A93FFFFFFFFFFDC9325DCB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hF5F5F5B5AC6C6464ADF6ADCA93DC0125258A014ADC9325254A4A932593DC1DDC),
    .INIT_1A(256'hABECF4F5F5F5B4ABA3A3ABECF5FEF5F5ECECECACF5F5FEF6F664932593921BF5),
    .INIT_1B(256'hE3A3AD65D325B664ACECECECECECECECF4F4F4F5F5F5F5F5F5F5F5F5F5ACAC63),
    .INIT_1C(256'h241B241BDA23FFFFB69365A3A3A3A4A464A4A3A3A35BD39494534A0012A3A3A3),
    .INIT_1D(256'hABA3ABECACACF4F5FEFEFEFDF5F5F5FEFEFEFEFEFEFEFDACF5FEF589DB9292DB),
    .INIT_1E(256'hFFFFFFFFFFFFF6F5F4A3ABAB1A63FEFEFDF5ABACFDFDF5F5FDF5F5F4ACACACEC),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_061440_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n116 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i60_008,inst_doa_i60_007,inst_doa_i60_006,inst_doa_i60_005,inst_doa_i60_004,inst_doa_i60_003,inst_doa_i60_002,inst_doa_i60_001,inst_doa_i60_000}));
  // address_offset=62464;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFE1F3BFFE0FF7FFFFFFFFFFFFC1FFF183123F5FFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFF1B71FFF1FFFFFFFFFFFFFFFE9FFF982123FAFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFF9B71FFFFFFBFFFFFFFFFFFFE0FFF982123FAFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFF1B71FFFFFFFFFFFFFFFFFFFE0FFF982121FCFFFFF),
    .INIT_00(256'h9300B6FFFFFFFFB68B25DC25FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFEFEFEFEFEFEFEB56464B5ADDCDC012525930093DC93251D4A4A932593DC25DC),
    .INIT_02(256'hACF4F5FEFEF5F5F4ABA3ABABACF5FEFEF5ACF5F6FEFEFEF5F5B592DCDC4A92B5),
    .INIT_03(256'hE3A36C24DC6E6E6DACECECECECECECF4F4F5F5F5F5F5F5F5F5F5F5F5F5ACACAC),
    .INIT_04(256'h24236C23DADBFFFF254A2464A3E3ECECEDECECECE3A31B4A535300D2A3A3A3A3),
    .INIT_05(256'hA3ABECACABECF5FEFEFEFEF5F5F5FDFEFEFEFEFEFFFEF5ACFDFEB500DB92DB1B),
    .INIT_06(256'hFFFFFFFFFFFFF5FDF5A3ABAB1A6CFEFEFDF5ABACFDFEFEF5FDF5F4F4ACABABAB),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h93006EFFFFFFFFFF259325DCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFEFEFEFEFEFEFEFEFEF56C6D6DDC012525930093DC9326DC4A4A932593DC25DC),
    .INIT_0A(256'hACF5F5FEFEFEFEFEFEF4ABABABECF5FDFEFEFEFFFFFEFEFEFDF5248A1D930165),
    .INIT_0B(256'hECAC6C656E2625B6ACECECECECECF4F4F5F5F5F5F6F5F5F5F5F5F5F5F5ECECAC),
    .INIT_0C(256'h24DB6D24D21BFFFF9393DC6DACECECECECECECECECECA41B920092A4ECECECEC),
    .INIT_0D(256'hA3ECABABACF5F5FEFEFEF5F4F5F5FEFEFEFEFEFEFFFEF5B5FEFEB564DB92DA23),
    .INIT_0E(256'hFFFFFFFFFFFFF5FDF5A3A3AB1A6CFEFDFDF5ACABF5FEFEFDF5F5F4F4ACABABA3),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hD30025FFFFFFFFFFB7931DDCB6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hF5FEFEFEFEFEFEFEFEFEFE6D6DD30125259301DCD49366DC4A4A932593DC25DC),
    .INIT_12(256'hACF5FDFEFEFEFEFEFEFEFDACABACACF5FDFEFEFEFEFEFEFEFEFEB549DCDC01DC),
    .INIT_13(256'hECF5ACAD6EDD6EADACECECECECF4F5F5F5F5F5F5F5F6F6F6F6F6F6F5F5ECACAC),
    .INIT_14(256'h24DBB624921BFFB6424BDCAEACECECECECECECECECECEDEDAC63ACEDEDF5ECF4),
    .INIT_15(256'hABECABABF4F5FDFEFDF5F5F4F5FDFEFEFEFEFEFEFFFEF5FDFEFEACB51B92DB23),
    .INIT_16(256'hFFFFFFFFFFFEF5F5F5ABA3AB1AACFEFDFDF5F4ABF5FDFEFDF5F5F4ECABABA3A3),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hD341DBFFFFFFFFFFFF25D4DD25FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hB4FEF5FEFEFEFEFEFEFEFEFE6D924A65254A4ADC93DC66934A8A932593DC25DC),
    .INIT_1A(256'hACF5FDFEFEFEFEFEFEFEFEF5ACACACECF5FDFEFEFEFEFEFEFEFEFE9293DD8B8A),
    .INIT_1B(256'hECF4ECAD65262524ACECECECECF4F4F5F5F5F5F5FEFEFEFEFEF6F5F5F5F5ECAC),
    .INIT_1C(256'h2492FF6D8923FF254A8BDC6DADECECECECECECECECEDEDF4F4F5F5F5F5F5F5F5),
    .INIT_1D(256'hECABABB4F5FDFDFDF5F4F4F5F5FEFEFEFEFEFEFEFEFEF5F5FEF5B4F5D292DB23),
    .INIT_1E(256'hFFFFFFFFFFFEF5F5F5ACA3AB63ACFEF5FDFDF4ABECF5FDFDF5F5ECACABA3A3A3),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_062464_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n116 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i61_008,inst_doa_i61_007,inst_doa_i61_006,inst_doa_i61_005,inst_doa_i61_004,inst_doa_i61_003,inst_doa_i61_002,inst_doa_i61_001,inst_doa_i61_000}));
  // address_offset=63488;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFF1B63FFFFFFDFFFFFFFFFFFFF0FFF986121FC7FFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFF1763FFFFFFCFFFFFFFFFFFFF0FFFD06121FC7FFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFF17627FFFFFCFFFFFFFFFFFFF07FFF04035FC7FFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFF96E27FFFFFCFFFFFFFFFFFFF07FFF04035FEBFFFF),
    .INIT_00(256'hD49392FFFFFFFFFFFFB693DDDCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h6CFDF5FDFEFEFEFEFEFEFEFEFEE34A6E1C4A93DC4A2525938A938A2593D425DC),
    .INIT_02(256'hACF5FDFEFEFEFEFEFEFEFEFEF5ACF4F4F4F5FDFEFEFEFEFEFEFEFE2401DCDC01),
    .INIT_03(256'hF5F4ECACAE6E931C64ECECECECF4F5F5F5F5F5FDFDFEFEFEFEF6F6F6F5F5ECAC),
    .INIT_04(256'h23DBFF64496CFFDC4B931D6565ACECECECECECECEDEDECF4F5F5F5F5F5F5F5F5),
    .INIT_05(256'hABABACF5FDFDFDF5F4F4F4F5FEFEFEFEFEFEFEFEFEF5ACFDFEACF5AC4892DB64),
    .INIT_06(256'hFFFFFFFFFFF6F5F5F5ECA3A363B4FDF5F5F5F5ACECF4F5FDF5F4ACABA3A362AB),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hDCDC4AB6FFFFFFFFFFF7DBDCDC6EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h23F5F5F5FDFEFEFEFEFEFEFEFEB6DC6EDC4AD4934B25259392938A1C93D425DD),
    .INIT_0A(256'hACF5FEFEFEFEFEFEFEFEFEFEFEFDACF4ECF4F5F5FDFEFEFEFEFEFF6D01DCDC01),
    .INIT_0B(256'hF5F5F5ECAD254BDB64ACECECECF5F5F5F5F5F6FEFEFEFEFEFEFEF6F6F6F5EDED),
    .INIT_0C(256'hDB2CFF2491B5B6935393251C2464ECECECECECECEDF5F5F5F5F5F5F5F5F5F5F5),
    .INIT_0D(256'hABACF4F5F5F5F5F4F4F4F5F5FEFEFEFEFEFEFEFEFEB4F4FEFEF5FDAC49DBDB6C),
    .INIT_0E(256'hFFFFFFFFFFF6F5F5F5F4A3A363B4FDF5F5F5F5ACF4ECF4F5F5ECACABA362ABAB),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h9325936DFFFFFFFFFFFFDCDCDD25FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hDAFEFEF5FDFEFDFEFEFEFEFEFEFF6D26DC93DC4A9466DC938A934ADC93D42525),
    .INIT_12(256'hACF5FEFEFEFEFEFEFEFEFEFEFEFEF5ACF4ECF4F5F5FDFEFEFEFEFF6D0194DC01),
    .INIT_13(256'hF5F5F5F5AC2493936DADECECEDF5F5F5F6F6FEFEFEFEFEFEFEFEFEF6F6F5F5ED),
    .INIT_14(256'hDB6DFF1BDAFE6E4A4BDC25DCDC64ACECECECECECF4F5F5F5F5F5F5F5F5F5F5F5),
    .INIT_15(256'hACF4F5FDF5F4F4F4F4F4F5FEFEFEFEFEFEFEFEFEFEACFDFEB5F5F5ACD2DBDB6C),
    .INIT_16(256'hFFFFFFFFFFF5F5F5F5F5AB62A3F4F5F4F5F5F5ACF4ACACF4F4ECABA3A262ACAB),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h9365DC6DFFFFFFFFFFFF244A1DDCF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h49BEFEFEFEFEFDFDFEFEFEFEFEFEF62493D3934ADC25DC938A934ADC93DC2525),
    .INIT_1A(256'hACF5FEFEFEFEFEFEFEFEFEFEF5FDFEF5ECF4ECF4F5F5FDFEFEFEFF6D0194D492),
    .INIT_1B(256'hF5F5F5F5AC6492DCB6ADECECEDF5F5F5F6F6FEFEFEFEFEFEFEFEFEF6F6F5F5F5),
    .INIT_1C(256'hDBFFFFDB24FF254A4BDC25D4931C64ACECECECECF4F4F5F5F5F5F5F5F5F5F5F5),
    .INIT_1D(256'hF4F5F5F5F4ECECF4F4F5FDFEFEFEFEFEFEFEFEFEF5B4FEF5F5FDF4AC2392DB24),
    .INIT_1E(256'hFFFFFFFFFEF5F5F5F5F5EC62A3F4F5F4F5F5F5B4F4ACACACF4ECABA3A3ABABAC),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_063488_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n116 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i62_008,inst_doa_i62_007,inst_doa_i62_006,inst_doa_i62_005,inst_doa_i62_004,inst_doa_i62_003,inst_doa_i62_002,inst_doa_i62_001,inst_doa_i62_000}));
  // address_offset=64512;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=9;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFBEC63FFFFFDFFFFFFFFFFFFF07FFF0C037FE3FFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFBEC41FFFFFF7FFFFFFFFFFFF07FFF08036FE3FFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFBEC41FFFFFE7FFFFFFFFFFFF07FFF08036FE1FFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFE840FFFFFE7FFFFFFFFFFFF07FFF98036FE1FFFF),
    .INIT_00(256'h936E2524FFFFFFFFFFFF6D00DCDC6EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h00B6FFFEFEFEFEFDFEFEFEFEFEFEFF6493DC4A932525DC9393934ADC4ADC2525),
    .INIT_02(256'hECF5FDFEFEFEFEFEFEFEFEFEFDF5F5FEF5F4F4F4F4F4F5FDFDFEFE6D0193D393),
    .INIT_03(256'hF5F5F5F5F564DC2E2564ECECEDF5F5F5F6F6FEFEFEFEFEFEFEFEFEFEF5F5F5F5),
    .INIT_04(256'h6DFFFFDB24BFDC4B93251D948B9324ACECECECECF4F4F5F5F5F5F5F5F6F6F6F5),
    .INIT_05(256'hF5F5F5F4ECECF4F4F4FDFEFEFEFEFEFEFEFEFEFEB5FDFEB5FEF5B4F564492324),
    .INIT_06(256'hFFFFFFFFFEF5F5F5F5F5F4A3A3F4F5F4F4F5F5F4F4ACACACACEBABA3A3ABABF4),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h8B6E6EDBFFFFFFFFFFFF6E0093DC24FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h00B6FFFEFEFEFEFEFEFEFEFEFEFEFEB593934ADC25DCDB9393934ADC4ADC2525),
    .INIT_0A(256'hF4F5FDFEFEFEFEFEFEFEFEFEFEF5B4FDFEF4F5F4ECF4F4F5F5F5FE6D01939393),
    .INIT_0B(256'hF5F5F5F5F5AD6D259324ACF4ECF5F5F5F6FEFEFEFEFEFEFEFEFEFEFEFDF5F5F5),
    .INIT_0C(256'hB6FFF7496DB6938B9325DC938B93DB64ECECECECF5F4F5F5F6F6F6F6FEFEF6F6),
    .INIT_0D(256'hF5F4F4ECECECECF4F5FEFEFEFEFEFEFEFEFEFEFEF5FEB5F5FEF5F5FEAD48242C),
    .INIT_0E(256'hFFFFFFFFF6F5F5F4F4F4F4ABA3F4F5F4F4F5F4F4F4AC6DADABABABA3ABABECF5),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h936EB692FFFFFFFFFFFFB64149DCDCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h006DFFFEFEFEFEFEFEFEFEFEFEFEFEFEDB0193DD26DCDC8A93934ADC4ADC2525),
    .INIT_12(256'hF4F5FDFEFEFEFEFEFEFEFEFEFEF5ACF4FDFEB4F5ECECF4F4F5F5FD64499493DB),
    .INIT_13(256'hF5F5F5F5F5EDAE934A24ACF4F4F5F5F5F6FEFEFEFEFEFEFEFEFEFEFEFEF5F5F5),
    .INIT_14(256'hFFFFB6492C6D934BD425DC939393921CACEDECECF4F4F5F5F6F6F6F6FEFEFEF6),
    .INIT_15(256'hF4ECACECF4ECF4F5FEFEFEFEFEFEFEFEFEFEFEF6FEFEB5FEFDFDFEFEFEDA246D),
    .INIT_16(256'hFFFFFFFFF5F5F5F4F4F4F4ACABF4F4B4F4F4F4F4F5AD6D6DABA2A3A3ECECF4F5),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h936EB749B7FFFFFFFFFFB78A00DBDC6EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h0025FFFEFEFEFEFEFEFEFEFEFEFEFEFF6E01DC2525DCDB4AD34A8BD34ADC2525),
    .INIT_1A(256'hF4F5FEFEFEFEFEFEFEFEFEFEFEFEF4ACB4FDF5ECF5ECECF4F4F5F52392944ADC),
    .INIT_1B(256'hFEF6F6F5F5F56D93931BA4F4F5F5F5F6FDFEFEFEFEFEFEFFFFFEFEFEFEF6F5F6),
    .INIT_1C(256'hFFFFB69224DC934ADC259352939201DC64ECF4F4F4F4F5F5F5F6F6F6FEFEFEFE),
    .INIT_1D(256'hACACECECECECF5FDFEFEFEFEFEFEFEFEFEFEFEF5FEF5FEFEFDFEFEFEFE6C6DB6),
    .INIT_1E(256'hFFFFFFFFF5F5F5F4F4F4F4ACABF4F4ACECF4B4F4F5AD656DA3A2A2ECECF4F4F4),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x9_sub_064512_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n116 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i63_008,inst_doa_i63_007,inst_doa_i63_006,inst_doa_i63_005,inst_doa_i63_004,inst_doa_i63_003,inst_doa_i63_002,inst_doa_i63_001,inst_doa_i63_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_10  (
    .i0(inst_doa_i20_000),
    .i1(inst_doa_i21_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_10 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_11  (
    .i0(inst_doa_i22_000),
    .i1(inst_doa_i23_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_11 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_12  (
    .i0(inst_doa_i24_000),
    .i1(inst_doa_i25_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_12 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_13  (
    .i0(inst_doa_i26_000),
    .i1(inst_doa_i27_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_13 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_14  (
    .i0(inst_doa_i28_000),
    .i1(inst_doa_i29_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_14 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_15  (
    .i0(inst_doa_i30_000),
    .i1(inst_doa_i31_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_15 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_16  (
    .i0(inst_doa_i32_000),
    .i1(inst_doa_i33_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_16 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_17  (
    .i0(inst_doa_i34_000),
    .i1(inst_doa_i35_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_17 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_18  (
    .i0(inst_doa_i36_000),
    .i1(inst_doa_i37_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_18 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_19  (
    .i0(inst_doa_i38_000),
    .i1(inst_doa_i39_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_19 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_2  (
    .i0(inst_doa_i4_000),
    .i1(inst_doa_i5_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_20  (
    .i0(inst_doa_i40_000),
    .i1(inst_doa_i41_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_20 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_21  (
    .i0(inst_doa_i42_000),
    .i1(inst_doa_i43_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_21 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_22  (
    .i0(inst_doa_i44_000),
    .i1(inst_doa_i45_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_22 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_23  (
    .i0(inst_doa_i46_000),
    .i1(inst_doa_i47_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_23 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_24  (
    .i0(inst_doa_i48_000),
    .i1(inst_doa_i49_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_24 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_25  (
    .i0(inst_doa_i50_000),
    .i1(inst_doa_i51_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_25 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_26  (
    .i0(inst_doa_i52_000),
    .i1(inst_doa_i53_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_26 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_27  (
    .i0(inst_doa_i54_000),
    .i1(inst_doa_i55_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_27 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_28  (
    .i0(inst_doa_i56_000),
    .i1(inst_doa_i57_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_28 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_29  (
    .i0(inst_doa_i58_000),
    .i1(inst_doa_i59_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_29 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_3  (
    .i0(inst_doa_i6_000),
    .i1(inst_doa_i7_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_30  (
    .i0(inst_doa_i60_000),
    .i1(inst_doa_i61_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_30 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_31  (
    .i0(inst_doa_i62_000),
    .i1(inst_doa_i63_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_31 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_4  (
    .i0(inst_doa_i8_000),
    .i1(inst_doa_i9_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_4 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_5  (
    .i0(inst_doa_i10_000),
    .i1(inst_doa_i11_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_5 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_6  (
    .i0(inst_doa_i12_000),
    .i1(inst_doa_i13_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_6 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_7  (
    .i0(inst_doa_i14_000),
    .i1(inst_doa_i15_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_7 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_8  (
    .i0(inst_doa_i16_000),
    .i1(inst_doa_i17_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_8 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_9  (
    .i0(inst_doa_i18_000),
    .i1(inst_doa_i19_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_9 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b0/B0_2 ),
    .i1(\inst_doa_mux_b0/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b0/B0_20 ),
    .i1(\inst_doa_mux_b0/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_10 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b0/B0_22 ),
    .i1(\inst_doa_mux_b0/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_11 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b0/B0_24 ),
    .i1(\inst_doa_mux_b0/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_12 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b0/B0_26 ),
    .i1(\inst_doa_mux_b0/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_13 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b0/B0_28 ),
    .i1(\inst_doa_mux_b0/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_14 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b0/B0_30 ),
    .i1(\inst_doa_mux_b0/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_15 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b0/B0_4 ),
    .i1(\inst_doa_mux_b0/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b0/B0_6 ),
    .i1(\inst_doa_mux_b0/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b0/B0_8 ),
    .i1(\inst_doa_mux_b0/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_4 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b0/B0_10 ),
    .i1(\inst_doa_mux_b0/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_5 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b0/B0_12 ),
    .i1(\inst_doa_mux_b0/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_6 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b0/B0_14 ),
    .i1(\inst_doa_mux_b0/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_7 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b0/B0_16 ),
    .i1(\inst_doa_mux_b0/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_8 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b0/B0_18 ),
    .i1(\inst_doa_mux_b0/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_9 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b0/B1_0 ),
    .i1(\inst_doa_mux_b0/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b0/B1_2 ),
    .i1(\inst_doa_mux_b0/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b0/B1_4 ),
    .i1(\inst_doa_mux_b0/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b0/B1_6 ),
    .i1(\inst_doa_mux_b0/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b0/B1_8 ),
    .i1(\inst_doa_mux_b0/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_4 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b0/B1_10 ),
    .i1(\inst_doa_mux_b0/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_5 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b0/B1_12 ),
    .i1(\inst_doa_mux_b0/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_6 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b0/B1_14 ),
    .i1(\inst_doa_mux_b0/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_7 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b0/B2_0 ),
    .i1(\inst_doa_mux_b0/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b0/B3_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b0/B2_2 ),
    .i1(\inst_doa_mux_b0/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b0/B3_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b0/B2_4 ),
    .i1(\inst_doa_mux_b0/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b0/B3_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b0/B2_6 ),
    .i1(\inst_doa_mux_b0/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b0/B3_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b0/B3_0 ),
    .i1(\inst_doa_mux_b0/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b0/B4_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b0/B3_2 ),
    .i1(\inst_doa_mux_b0/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b0/B4_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b0/B4_0 ),
    .i1(\inst_doa_mux_b0/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_10  (
    .i0(inst_doa_i20_001),
    .i1(inst_doa_i21_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_10 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_11  (
    .i0(inst_doa_i22_001),
    .i1(inst_doa_i23_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_11 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_12  (
    .i0(inst_doa_i24_001),
    .i1(inst_doa_i25_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_12 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_13  (
    .i0(inst_doa_i26_001),
    .i1(inst_doa_i27_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_13 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_14  (
    .i0(inst_doa_i28_001),
    .i1(inst_doa_i29_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_14 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_15  (
    .i0(inst_doa_i30_001),
    .i1(inst_doa_i31_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_15 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_16  (
    .i0(inst_doa_i32_001),
    .i1(inst_doa_i33_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_16 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_17  (
    .i0(inst_doa_i34_001),
    .i1(inst_doa_i35_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_17 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_18  (
    .i0(inst_doa_i36_001),
    .i1(inst_doa_i37_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_18 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_19  (
    .i0(inst_doa_i38_001),
    .i1(inst_doa_i39_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_19 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_2  (
    .i0(inst_doa_i4_001),
    .i1(inst_doa_i5_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_20  (
    .i0(inst_doa_i40_001),
    .i1(inst_doa_i41_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_20 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_21  (
    .i0(inst_doa_i42_001),
    .i1(inst_doa_i43_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_21 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_22  (
    .i0(inst_doa_i44_001),
    .i1(inst_doa_i45_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_22 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_23  (
    .i0(inst_doa_i46_001),
    .i1(inst_doa_i47_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_23 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_24  (
    .i0(inst_doa_i48_001),
    .i1(inst_doa_i49_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_24 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_25  (
    .i0(inst_doa_i50_001),
    .i1(inst_doa_i51_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_25 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_26  (
    .i0(inst_doa_i52_001),
    .i1(inst_doa_i53_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_26 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_27  (
    .i0(inst_doa_i54_001),
    .i1(inst_doa_i55_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_27 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_28  (
    .i0(inst_doa_i56_001),
    .i1(inst_doa_i57_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_28 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_29  (
    .i0(inst_doa_i58_001),
    .i1(inst_doa_i59_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_29 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_3  (
    .i0(inst_doa_i6_001),
    .i1(inst_doa_i7_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_30  (
    .i0(inst_doa_i60_001),
    .i1(inst_doa_i61_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_30 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_31  (
    .i0(inst_doa_i62_001),
    .i1(inst_doa_i63_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_31 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_4  (
    .i0(inst_doa_i8_001),
    .i1(inst_doa_i9_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_4 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_5  (
    .i0(inst_doa_i10_001),
    .i1(inst_doa_i11_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_5 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_6  (
    .i0(inst_doa_i12_001),
    .i1(inst_doa_i13_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_6 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_7  (
    .i0(inst_doa_i14_001),
    .i1(inst_doa_i15_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_7 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_8  (
    .i0(inst_doa_i16_001),
    .i1(inst_doa_i17_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_8 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_9  (
    .i0(inst_doa_i18_001),
    .i1(inst_doa_i19_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_9 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b1/B0_2 ),
    .i1(\inst_doa_mux_b1/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b1/B0_20 ),
    .i1(\inst_doa_mux_b1/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_10 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b1/B0_22 ),
    .i1(\inst_doa_mux_b1/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_11 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b1/B0_24 ),
    .i1(\inst_doa_mux_b1/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_12 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b1/B0_26 ),
    .i1(\inst_doa_mux_b1/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_13 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b1/B0_28 ),
    .i1(\inst_doa_mux_b1/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_14 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b1/B0_30 ),
    .i1(\inst_doa_mux_b1/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_15 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b1/B0_4 ),
    .i1(\inst_doa_mux_b1/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b1/B0_6 ),
    .i1(\inst_doa_mux_b1/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b1/B0_8 ),
    .i1(\inst_doa_mux_b1/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_4 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b1/B0_10 ),
    .i1(\inst_doa_mux_b1/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_5 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b1/B0_12 ),
    .i1(\inst_doa_mux_b1/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_6 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b1/B0_14 ),
    .i1(\inst_doa_mux_b1/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_7 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b1/B0_16 ),
    .i1(\inst_doa_mux_b1/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_8 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b1/B0_18 ),
    .i1(\inst_doa_mux_b1/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_9 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b1/B1_0 ),
    .i1(\inst_doa_mux_b1/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b1/B1_2 ),
    .i1(\inst_doa_mux_b1/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b1/B1_4 ),
    .i1(\inst_doa_mux_b1/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b1/B1_6 ),
    .i1(\inst_doa_mux_b1/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b1/B1_8 ),
    .i1(\inst_doa_mux_b1/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_4 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b1/B1_10 ),
    .i1(\inst_doa_mux_b1/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_5 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b1/B1_12 ),
    .i1(\inst_doa_mux_b1/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_6 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b1/B1_14 ),
    .i1(\inst_doa_mux_b1/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_7 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b1/B2_0 ),
    .i1(\inst_doa_mux_b1/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b1/B3_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b1/B2_2 ),
    .i1(\inst_doa_mux_b1/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b1/B3_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b1/B2_4 ),
    .i1(\inst_doa_mux_b1/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b1/B3_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b1/B2_6 ),
    .i1(\inst_doa_mux_b1/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b1/B3_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b1/B3_0 ),
    .i1(\inst_doa_mux_b1/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b1/B4_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b1/B3_2 ),
    .i1(\inst_doa_mux_b1/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b1/B4_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b1/B4_0 ),
    .i1(\inst_doa_mux_b1/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_10  (
    .i0(inst_doa_i20_002),
    .i1(inst_doa_i21_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_10 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_11  (
    .i0(inst_doa_i22_002),
    .i1(inst_doa_i23_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_11 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_12  (
    .i0(inst_doa_i24_002),
    .i1(inst_doa_i25_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_12 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_13  (
    .i0(inst_doa_i26_002),
    .i1(inst_doa_i27_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_13 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_14  (
    .i0(inst_doa_i28_002),
    .i1(inst_doa_i29_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_14 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_15  (
    .i0(inst_doa_i30_002),
    .i1(inst_doa_i31_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_15 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_16  (
    .i0(inst_doa_i32_002),
    .i1(inst_doa_i33_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_16 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_17  (
    .i0(inst_doa_i34_002),
    .i1(inst_doa_i35_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_17 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_18  (
    .i0(inst_doa_i36_002),
    .i1(inst_doa_i37_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_18 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_19  (
    .i0(inst_doa_i38_002),
    .i1(inst_doa_i39_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_19 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_2  (
    .i0(inst_doa_i4_002),
    .i1(inst_doa_i5_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_20  (
    .i0(inst_doa_i40_002),
    .i1(inst_doa_i41_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_20 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_21  (
    .i0(inst_doa_i42_002),
    .i1(inst_doa_i43_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_21 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_22  (
    .i0(inst_doa_i44_002),
    .i1(inst_doa_i45_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_22 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_23  (
    .i0(inst_doa_i46_002),
    .i1(inst_doa_i47_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_23 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_24  (
    .i0(inst_doa_i48_002),
    .i1(inst_doa_i49_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_24 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_25  (
    .i0(inst_doa_i50_002),
    .i1(inst_doa_i51_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_25 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_26  (
    .i0(inst_doa_i52_002),
    .i1(inst_doa_i53_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_26 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_27  (
    .i0(inst_doa_i54_002),
    .i1(inst_doa_i55_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_27 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_28  (
    .i0(inst_doa_i56_002),
    .i1(inst_doa_i57_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_28 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_29  (
    .i0(inst_doa_i58_002),
    .i1(inst_doa_i59_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_29 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_3  (
    .i0(inst_doa_i6_002),
    .i1(inst_doa_i7_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_30  (
    .i0(inst_doa_i60_002),
    .i1(inst_doa_i61_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_30 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_31  (
    .i0(inst_doa_i62_002),
    .i1(inst_doa_i63_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_31 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_4  (
    .i0(inst_doa_i8_002),
    .i1(inst_doa_i9_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_4 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_5  (
    .i0(inst_doa_i10_002),
    .i1(inst_doa_i11_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_5 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_6  (
    .i0(inst_doa_i12_002),
    .i1(inst_doa_i13_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_6 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_7  (
    .i0(inst_doa_i14_002),
    .i1(inst_doa_i15_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_7 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_8  (
    .i0(inst_doa_i16_002),
    .i1(inst_doa_i17_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_8 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_9  (
    .i0(inst_doa_i18_002),
    .i1(inst_doa_i19_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_9 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b2/B0_2 ),
    .i1(\inst_doa_mux_b2/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b2/B0_20 ),
    .i1(\inst_doa_mux_b2/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_10 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b2/B0_22 ),
    .i1(\inst_doa_mux_b2/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_11 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b2/B0_24 ),
    .i1(\inst_doa_mux_b2/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_12 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b2/B0_26 ),
    .i1(\inst_doa_mux_b2/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_13 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b2/B0_28 ),
    .i1(\inst_doa_mux_b2/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_14 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b2/B0_30 ),
    .i1(\inst_doa_mux_b2/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_15 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b2/B0_4 ),
    .i1(\inst_doa_mux_b2/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b2/B0_6 ),
    .i1(\inst_doa_mux_b2/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b2/B0_8 ),
    .i1(\inst_doa_mux_b2/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_4 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b2/B0_10 ),
    .i1(\inst_doa_mux_b2/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_5 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b2/B0_12 ),
    .i1(\inst_doa_mux_b2/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_6 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b2/B0_14 ),
    .i1(\inst_doa_mux_b2/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_7 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b2/B0_16 ),
    .i1(\inst_doa_mux_b2/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_8 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b2/B0_18 ),
    .i1(\inst_doa_mux_b2/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_9 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b2/B1_0 ),
    .i1(\inst_doa_mux_b2/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b2/B1_2 ),
    .i1(\inst_doa_mux_b2/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b2/B1_4 ),
    .i1(\inst_doa_mux_b2/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b2/B1_6 ),
    .i1(\inst_doa_mux_b2/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b2/B1_8 ),
    .i1(\inst_doa_mux_b2/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_4 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b2/B1_10 ),
    .i1(\inst_doa_mux_b2/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_5 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b2/B1_12 ),
    .i1(\inst_doa_mux_b2/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_6 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b2/B1_14 ),
    .i1(\inst_doa_mux_b2/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_7 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b2/B2_0 ),
    .i1(\inst_doa_mux_b2/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b2/B3_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b2/B2_2 ),
    .i1(\inst_doa_mux_b2/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b2/B3_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b2/B2_4 ),
    .i1(\inst_doa_mux_b2/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b2/B3_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b2/B2_6 ),
    .i1(\inst_doa_mux_b2/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b2/B3_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b2/B3_0 ),
    .i1(\inst_doa_mux_b2/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b2/B4_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b2/B3_2 ),
    .i1(\inst_doa_mux_b2/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b2/B4_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b2/B4_0 ),
    .i1(\inst_doa_mux_b2/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_10  (
    .i0(inst_doa_i20_003),
    .i1(inst_doa_i21_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_10 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_11  (
    .i0(inst_doa_i22_003),
    .i1(inst_doa_i23_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_11 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_12  (
    .i0(inst_doa_i24_003),
    .i1(inst_doa_i25_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_12 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_13  (
    .i0(inst_doa_i26_003),
    .i1(inst_doa_i27_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_13 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_14  (
    .i0(inst_doa_i28_003),
    .i1(inst_doa_i29_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_14 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_15  (
    .i0(inst_doa_i30_003),
    .i1(inst_doa_i31_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_15 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_16  (
    .i0(inst_doa_i32_003),
    .i1(inst_doa_i33_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_16 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_17  (
    .i0(inst_doa_i34_003),
    .i1(inst_doa_i35_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_17 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_18  (
    .i0(inst_doa_i36_003),
    .i1(inst_doa_i37_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_18 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_19  (
    .i0(inst_doa_i38_003),
    .i1(inst_doa_i39_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_19 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_2  (
    .i0(inst_doa_i4_003),
    .i1(inst_doa_i5_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_2 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_20  (
    .i0(inst_doa_i40_003),
    .i1(inst_doa_i41_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_20 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_21  (
    .i0(inst_doa_i42_003),
    .i1(inst_doa_i43_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_21 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_22  (
    .i0(inst_doa_i44_003),
    .i1(inst_doa_i45_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_22 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_23  (
    .i0(inst_doa_i46_003),
    .i1(inst_doa_i47_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_23 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_24  (
    .i0(inst_doa_i48_003),
    .i1(inst_doa_i49_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_24 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_25  (
    .i0(inst_doa_i50_003),
    .i1(inst_doa_i51_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_25 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_26  (
    .i0(inst_doa_i52_003),
    .i1(inst_doa_i53_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_26 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_27  (
    .i0(inst_doa_i54_003),
    .i1(inst_doa_i55_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_27 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_28  (
    .i0(inst_doa_i56_003),
    .i1(inst_doa_i57_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_28 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_29  (
    .i0(inst_doa_i58_003),
    .i1(inst_doa_i59_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_29 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_3  (
    .i0(inst_doa_i6_003),
    .i1(inst_doa_i7_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_3 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_30  (
    .i0(inst_doa_i60_003),
    .i1(inst_doa_i61_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_30 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_31  (
    .i0(inst_doa_i62_003),
    .i1(inst_doa_i63_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_31 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_4  (
    .i0(inst_doa_i8_003),
    .i1(inst_doa_i9_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_4 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_5  (
    .i0(inst_doa_i10_003),
    .i1(inst_doa_i11_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_5 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_6  (
    .i0(inst_doa_i12_003),
    .i1(inst_doa_i13_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_6 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_7  (
    .i0(inst_doa_i14_003),
    .i1(inst_doa_i15_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_7 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_8  (
    .i0(inst_doa_i16_003),
    .i1(inst_doa_i17_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_8 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_9  (
    .i0(inst_doa_i18_003),
    .i1(inst_doa_i19_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_9 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b3/B0_2 ),
    .i1(\inst_doa_mux_b3/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b3/B0_20 ),
    .i1(\inst_doa_mux_b3/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_10 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b3/B0_22 ),
    .i1(\inst_doa_mux_b3/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_11 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b3/B0_24 ),
    .i1(\inst_doa_mux_b3/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_12 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b3/B0_26 ),
    .i1(\inst_doa_mux_b3/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_13 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b3/B0_28 ),
    .i1(\inst_doa_mux_b3/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_14 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b3/B0_30 ),
    .i1(\inst_doa_mux_b3/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_15 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b3/B0_4 ),
    .i1(\inst_doa_mux_b3/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_2 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b3/B0_6 ),
    .i1(\inst_doa_mux_b3/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_3 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b3/B0_8 ),
    .i1(\inst_doa_mux_b3/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_4 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b3/B0_10 ),
    .i1(\inst_doa_mux_b3/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_5 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b3/B0_12 ),
    .i1(\inst_doa_mux_b3/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_6 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b3/B0_14 ),
    .i1(\inst_doa_mux_b3/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_7 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b3/B0_16 ),
    .i1(\inst_doa_mux_b3/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_8 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b3/B0_18 ),
    .i1(\inst_doa_mux_b3/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_9 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b3/B1_0 ),
    .i1(\inst_doa_mux_b3/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b3/B1_2 ),
    .i1(\inst_doa_mux_b3/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b3/B1_4 ),
    .i1(\inst_doa_mux_b3/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_2 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b3/B1_6 ),
    .i1(\inst_doa_mux_b3/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_3 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b3/B1_8 ),
    .i1(\inst_doa_mux_b3/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_4 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b3/B1_10 ),
    .i1(\inst_doa_mux_b3/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_5 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b3/B1_12 ),
    .i1(\inst_doa_mux_b3/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_6 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b3/B1_14 ),
    .i1(\inst_doa_mux_b3/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_7 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b3/B2_0 ),
    .i1(\inst_doa_mux_b3/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b3/B3_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b3/B2_2 ),
    .i1(\inst_doa_mux_b3/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b3/B3_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b3/B2_4 ),
    .i1(\inst_doa_mux_b3/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b3/B3_2 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b3/B2_6 ),
    .i1(\inst_doa_mux_b3/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b3/B3_3 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b3/B3_0 ),
    .i1(\inst_doa_mux_b3/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b3/B4_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b3/B3_2 ),
    .i1(\inst_doa_mux_b3/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b3/B4_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b3/B4_0 ),
    .i1(\inst_doa_mux_b3/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_10  (
    .i0(inst_doa_i20_004),
    .i1(inst_doa_i21_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_10 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_11  (
    .i0(inst_doa_i22_004),
    .i1(inst_doa_i23_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_11 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_12  (
    .i0(inst_doa_i24_004),
    .i1(inst_doa_i25_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_12 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_13  (
    .i0(inst_doa_i26_004),
    .i1(inst_doa_i27_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_13 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_14  (
    .i0(inst_doa_i28_004),
    .i1(inst_doa_i29_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_14 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_15  (
    .i0(inst_doa_i30_004),
    .i1(inst_doa_i31_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_15 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_16  (
    .i0(inst_doa_i32_004),
    .i1(inst_doa_i33_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_16 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_17  (
    .i0(inst_doa_i34_004),
    .i1(inst_doa_i35_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_17 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_18  (
    .i0(inst_doa_i36_004),
    .i1(inst_doa_i37_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_18 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_19  (
    .i0(inst_doa_i38_004),
    .i1(inst_doa_i39_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_19 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_2  (
    .i0(inst_doa_i4_004),
    .i1(inst_doa_i5_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_2 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_20  (
    .i0(inst_doa_i40_004),
    .i1(inst_doa_i41_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_20 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_21  (
    .i0(inst_doa_i42_004),
    .i1(inst_doa_i43_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_21 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_22  (
    .i0(inst_doa_i44_004),
    .i1(inst_doa_i45_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_22 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_23  (
    .i0(inst_doa_i46_004),
    .i1(inst_doa_i47_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_23 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_24  (
    .i0(inst_doa_i48_004),
    .i1(inst_doa_i49_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_24 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_25  (
    .i0(inst_doa_i50_004),
    .i1(inst_doa_i51_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_25 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_26  (
    .i0(inst_doa_i52_004),
    .i1(inst_doa_i53_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_26 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_27  (
    .i0(inst_doa_i54_004),
    .i1(inst_doa_i55_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_27 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_28  (
    .i0(inst_doa_i56_004),
    .i1(inst_doa_i57_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_28 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_29  (
    .i0(inst_doa_i58_004),
    .i1(inst_doa_i59_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_29 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_3  (
    .i0(inst_doa_i6_004),
    .i1(inst_doa_i7_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_3 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_30  (
    .i0(inst_doa_i60_004),
    .i1(inst_doa_i61_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_30 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_31  (
    .i0(inst_doa_i62_004),
    .i1(inst_doa_i63_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_31 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_4  (
    .i0(inst_doa_i8_004),
    .i1(inst_doa_i9_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_4 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_5  (
    .i0(inst_doa_i10_004),
    .i1(inst_doa_i11_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_5 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_6  (
    .i0(inst_doa_i12_004),
    .i1(inst_doa_i13_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_6 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_7  (
    .i0(inst_doa_i14_004),
    .i1(inst_doa_i15_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_7 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_8  (
    .i0(inst_doa_i16_004),
    .i1(inst_doa_i17_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_8 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_9  (
    .i0(inst_doa_i18_004),
    .i1(inst_doa_i19_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_9 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b4/B0_2 ),
    .i1(\inst_doa_mux_b4/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b4/B0_20 ),
    .i1(\inst_doa_mux_b4/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_10 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b4/B0_22 ),
    .i1(\inst_doa_mux_b4/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_11 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b4/B0_24 ),
    .i1(\inst_doa_mux_b4/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_12 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b4/B0_26 ),
    .i1(\inst_doa_mux_b4/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_13 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b4/B0_28 ),
    .i1(\inst_doa_mux_b4/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_14 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b4/B0_30 ),
    .i1(\inst_doa_mux_b4/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_15 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b4/B0_4 ),
    .i1(\inst_doa_mux_b4/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_2 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b4/B0_6 ),
    .i1(\inst_doa_mux_b4/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_3 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b4/B0_8 ),
    .i1(\inst_doa_mux_b4/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_4 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b4/B0_10 ),
    .i1(\inst_doa_mux_b4/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_5 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b4/B0_12 ),
    .i1(\inst_doa_mux_b4/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_6 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b4/B0_14 ),
    .i1(\inst_doa_mux_b4/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_7 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b4/B0_16 ),
    .i1(\inst_doa_mux_b4/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_8 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b4/B0_18 ),
    .i1(\inst_doa_mux_b4/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_9 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b4/B1_0 ),
    .i1(\inst_doa_mux_b4/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b4/B1_2 ),
    .i1(\inst_doa_mux_b4/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b4/B1_4 ),
    .i1(\inst_doa_mux_b4/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_2 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b4/B1_6 ),
    .i1(\inst_doa_mux_b4/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_3 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b4/B1_8 ),
    .i1(\inst_doa_mux_b4/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_4 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b4/B1_10 ),
    .i1(\inst_doa_mux_b4/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_5 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b4/B1_12 ),
    .i1(\inst_doa_mux_b4/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_6 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b4/B1_14 ),
    .i1(\inst_doa_mux_b4/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_7 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b4/B2_0 ),
    .i1(\inst_doa_mux_b4/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b4/B3_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b4/B2_2 ),
    .i1(\inst_doa_mux_b4/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b4/B3_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b4/B2_4 ),
    .i1(\inst_doa_mux_b4/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b4/B3_2 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b4/B2_6 ),
    .i1(\inst_doa_mux_b4/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b4/B3_3 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b4/B3_0 ),
    .i1(\inst_doa_mux_b4/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b4/B4_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b4/B3_2 ),
    .i1(\inst_doa_mux_b4/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b4/B4_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b4/B4_0 ),
    .i1(\inst_doa_mux_b4/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_10  (
    .i0(inst_doa_i20_005),
    .i1(inst_doa_i21_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_10 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_11  (
    .i0(inst_doa_i22_005),
    .i1(inst_doa_i23_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_11 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_12  (
    .i0(inst_doa_i24_005),
    .i1(inst_doa_i25_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_12 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_13  (
    .i0(inst_doa_i26_005),
    .i1(inst_doa_i27_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_13 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_14  (
    .i0(inst_doa_i28_005),
    .i1(inst_doa_i29_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_14 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_15  (
    .i0(inst_doa_i30_005),
    .i1(inst_doa_i31_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_15 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_16  (
    .i0(inst_doa_i32_005),
    .i1(inst_doa_i33_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_16 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_17  (
    .i0(inst_doa_i34_005),
    .i1(inst_doa_i35_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_17 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_18  (
    .i0(inst_doa_i36_005),
    .i1(inst_doa_i37_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_18 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_19  (
    .i0(inst_doa_i38_005),
    .i1(inst_doa_i39_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_19 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_2  (
    .i0(inst_doa_i4_005),
    .i1(inst_doa_i5_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_2 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_20  (
    .i0(inst_doa_i40_005),
    .i1(inst_doa_i41_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_20 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_21  (
    .i0(inst_doa_i42_005),
    .i1(inst_doa_i43_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_21 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_22  (
    .i0(inst_doa_i44_005),
    .i1(inst_doa_i45_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_22 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_23  (
    .i0(inst_doa_i46_005),
    .i1(inst_doa_i47_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_23 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_24  (
    .i0(inst_doa_i48_005),
    .i1(inst_doa_i49_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_24 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_25  (
    .i0(inst_doa_i50_005),
    .i1(inst_doa_i51_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_25 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_26  (
    .i0(inst_doa_i52_005),
    .i1(inst_doa_i53_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_26 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_27  (
    .i0(inst_doa_i54_005),
    .i1(inst_doa_i55_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_27 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_28  (
    .i0(inst_doa_i56_005),
    .i1(inst_doa_i57_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_28 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_29  (
    .i0(inst_doa_i58_005),
    .i1(inst_doa_i59_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_29 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_3  (
    .i0(inst_doa_i6_005),
    .i1(inst_doa_i7_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_3 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_30  (
    .i0(inst_doa_i60_005),
    .i1(inst_doa_i61_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_30 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_31  (
    .i0(inst_doa_i62_005),
    .i1(inst_doa_i63_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_31 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_4  (
    .i0(inst_doa_i8_005),
    .i1(inst_doa_i9_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_4 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_5  (
    .i0(inst_doa_i10_005),
    .i1(inst_doa_i11_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_5 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_6  (
    .i0(inst_doa_i12_005),
    .i1(inst_doa_i13_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_6 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_7  (
    .i0(inst_doa_i14_005),
    .i1(inst_doa_i15_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_7 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_8  (
    .i0(inst_doa_i16_005),
    .i1(inst_doa_i17_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_8 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_9  (
    .i0(inst_doa_i18_005),
    .i1(inst_doa_i19_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_9 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b5/B0_2 ),
    .i1(\inst_doa_mux_b5/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b5/B0_20 ),
    .i1(\inst_doa_mux_b5/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_10 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b5/B0_22 ),
    .i1(\inst_doa_mux_b5/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_11 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b5/B0_24 ),
    .i1(\inst_doa_mux_b5/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_12 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b5/B0_26 ),
    .i1(\inst_doa_mux_b5/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_13 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b5/B0_28 ),
    .i1(\inst_doa_mux_b5/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_14 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b5/B0_30 ),
    .i1(\inst_doa_mux_b5/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_15 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b5/B0_4 ),
    .i1(\inst_doa_mux_b5/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_2 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b5/B0_6 ),
    .i1(\inst_doa_mux_b5/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_3 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b5/B0_8 ),
    .i1(\inst_doa_mux_b5/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_4 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b5/B0_10 ),
    .i1(\inst_doa_mux_b5/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_5 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b5/B0_12 ),
    .i1(\inst_doa_mux_b5/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_6 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b5/B0_14 ),
    .i1(\inst_doa_mux_b5/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_7 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b5/B0_16 ),
    .i1(\inst_doa_mux_b5/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_8 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b5/B0_18 ),
    .i1(\inst_doa_mux_b5/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_9 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b5/B1_0 ),
    .i1(\inst_doa_mux_b5/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b5/B1_2 ),
    .i1(\inst_doa_mux_b5/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b5/B1_4 ),
    .i1(\inst_doa_mux_b5/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_2 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b5/B1_6 ),
    .i1(\inst_doa_mux_b5/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_3 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b5/B1_8 ),
    .i1(\inst_doa_mux_b5/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_4 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b5/B1_10 ),
    .i1(\inst_doa_mux_b5/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_5 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b5/B1_12 ),
    .i1(\inst_doa_mux_b5/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_6 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b5/B1_14 ),
    .i1(\inst_doa_mux_b5/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_7 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b5/B2_0 ),
    .i1(\inst_doa_mux_b5/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b5/B3_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b5/B2_2 ),
    .i1(\inst_doa_mux_b5/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b5/B3_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b5/B2_4 ),
    .i1(\inst_doa_mux_b5/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b5/B3_2 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b5/B2_6 ),
    .i1(\inst_doa_mux_b5/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b5/B3_3 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b5/B3_0 ),
    .i1(\inst_doa_mux_b5/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b5/B4_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b5/B3_2 ),
    .i1(\inst_doa_mux_b5/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b5/B4_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b5/B4_0 ),
    .i1(\inst_doa_mux_b5/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_10  (
    .i0(inst_doa_i20_006),
    .i1(inst_doa_i21_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_10 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_11  (
    .i0(inst_doa_i22_006),
    .i1(inst_doa_i23_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_11 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_12  (
    .i0(inst_doa_i24_006),
    .i1(inst_doa_i25_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_12 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_13  (
    .i0(inst_doa_i26_006),
    .i1(inst_doa_i27_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_13 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_14  (
    .i0(inst_doa_i28_006),
    .i1(inst_doa_i29_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_14 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_15  (
    .i0(inst_doa_i30_006),
    .i1(inst_doa_i31_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_15 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_16  (
    .i0(inst_doa_i32_006),
    .i1(inst_doa_i33_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_16 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_17  (
    .i0(inst_doa_i34_006),
    .i1(inst_doa_i35_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_17 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_18  (
    .i0(inst_doa_i36_006),
    .i1(inst_doa_i37_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_18 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_19  (
    .i0(inst_doa_i38_006),
    .i1(inst_doa_i39_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_19 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_2  (
    .i0(inst_doa_i4_006),
    .i1(inst_doa_i5_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_2 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_20  (
    .i0(inst_doa_i40_006),
    .i1(inst_doa_i41_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_20 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_21  (
    .i0(inst_doa_i42_006),
    .i1(inst_doa_i43_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_21 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_22  (
    .i0(inst_doa_i44_006),
    .i1(inst_doa_i45_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_22 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_23  (
    .i0(inst_doa_i46_006),
    .i1(inst_doa_i47_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_23 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_24  (
    .i0(inst_doa_i48_006),
    .i1(inst_doa_i49_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_24 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_25  (
    .i0(inst_doa_i50_006),
    .i1(inst_doa_i51_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_25 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_26  (
    .i0(inst_doa_i52_006),
    .i1(inst_doa_i53_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_26 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_27  (
    .i0(inst_doa_i54_006),
    .i1(inst_doa_i55_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_27 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_28  (
    .i0(inst_doa_i56_006),
    .i1(inst_doa_i57_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_28 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_29  (
    .i0(inst_doa_i58_006),
    .i1(inst_doa_i59_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_29 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_3  (
    .i0(inst_doa_i6_006),
    .i1(inst_doa_i7_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_3 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_30  (
    .i0(inst_doa_i60_006),
    .i1(inst_doa_i61_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_30 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_31  (
    .i0(inst_doa_i62_006),
    .i1(inst_doa_i63_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_31 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_4  (
    .i0(inst_doa_i8_006),
    .i1(inst_doa_i9_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_4 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_5  (
    .i0(inst_doa_i10_006),
    .i1(inst_doa_i11_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_5 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_6  (
    .i0(inst_doa_i12_006),
    .i1(inst_doa_i13_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_6 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_7  (
    .i0(inst_doa_i14_006),
    .i1(inst_doa_i15_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_7 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_8  (
    .i0(inst_doa_i16_006),
    .i1(inst_doa_i17_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_8 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_9  (
    .i0(inst_doa_i18_006),
    .i1(inst_doa_i19_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_9 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b6/B0_2 ),
    .i1(\inst_doa_mux_b6/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b6/B0_20 ),
    .i1(\inst_doa_mux_b6/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_10 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b6/B0_22 ),
    .i1(\inst_doa_mux_b6/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_11 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b6/B0_24 ),
    .i1(\inst_doa_mux_b6/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_12 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b6/B0_26 ),
    .i1(\inst_doa_mux_b6/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_13 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b6/B0_28 ),
    .i1(\inst_doa_mux_b6/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_14 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b6/B0_30 ),
    .i1(\inst_doa_mux_b6/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_15 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b6/B0_4 ),
    .i1(\inst_doa_mux_b6/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_2 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b6/B0_6 ),
    .i1(\inst_doa_mux_b6/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_3 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b6/B0_8 ),
    .i1(\inst_doa_mux_b6/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_4 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b6/B0_10 ),
    .i1(\inst_doa_mux_b6/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_5 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b6/B0_12 ),
    .i1(\inst_doa_mux_b6/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_6 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b6/B0_14 ),
    .i1(\inst_doa_mux_b6/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_7 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b6/B0_16 ),
    .i1(\inst_doa_mux_b6/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_8 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b6/B0_18 ),
    .i1(\inst_doa_mux_b6/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_9 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b6/B1_0 ),
    .i1(\inst_doa_mux_b6/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b6/B1_2 ),
    .i1(\inst_doa_mux_b6/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b6/B1_4 ),
    .i1(\inst_doa_mux_b6/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_2 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b6/B1_6 ),
    .i1(\inst_doa_mux_b6/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_3 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b6/B1_8 ),
    .i1(\inst_doa_mux_b6/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_4 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b6/B1_10 ),
    .i1(\inst_doa_mux_b6/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_5 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b6/B1_12 ),
    .i1(\inst_doa_mux_b6/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_6 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b6/B1_14 ),
    .i1(\inst_doa_mux_b6/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_7 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b6/B2_0 ),
    .i1(\inst_doa_mux_b6/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b6/B3_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b6/B2_2 ),
    .i1(\inst_doa_mux_b6/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b6/B3_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b6/B2_4 ),
    .i1(\inst_doa_mux_b6/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b6/B3_2 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b6/B2_6 ),
    .i1(\inst_doa_mux_b6/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b6/B3_3 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b6/B3_0 ),
    .i1(\inst_doa_mux_b6/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b6/B4_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b6/B3_2 ),
    .i1(\inst_doa_mux_b6/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b6/B4_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b6/B4_0 ),
    .i1(\inst_doa_mux_b6/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_10  (
    .i0(inst_doa_i20_007),
    .i1(inst_doa_i21_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_10 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_11  (
    .i0(inst_doa_i22_007),
    .i1(inst_doa_i23_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_11 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_12  (
    .i0(inst_doa_i24_007),
    .i1(inst_doa_i25_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_12 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_13  (
    .i0(inst_doa_i26_007),
    .i1(inst_doa_i27_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_13 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_14  (
    .i0(inst_doa_i28_007),
    .i1(inst_doa_i29_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_14 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_15  (
    .i0(inst_doa_i30_007),
    .i1(inst_doa_i31_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_15 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_16  (
    .i0(inst_doa_i32_007),
    .i1(inst_doa_i33_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_16 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_17  (
    .i0(inst_doa_i34_007),
    .i1(inst_doa_i35_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_17 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_18  (
    .i0(inst_doa_i36_007),
    .i1(inst_doa_i37_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_18 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_19  (
    .i0(inst_doa_i38_007),
    .i1(inst_doa_i39_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_19 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_2  (
    .i0(inst_doa_i4_007),
    .i1(inst_doa_i5_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_2 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_20  (
    .i0(inst_doa_i40_007),
    .i1(inst_doa_i41_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_20 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_21  (
    .i0(inst_doa_i42_007),
    .i1(inst_doa_i43_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_21 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_22  (
    .i0(inst_doa_i44_007),
    .i1(inst_doa_i45_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_22 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_23  (
    .i0(inst_doa_i46_007),
    .i1(inst_doa_i47_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_23 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_24  (
    .i0(inst_doa_i48_007),
    .i1(inst_doa_i49_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_24 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_25  (
    .i0(inst_doa_i50_007),
    .i1(inst_doa_i51_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_25 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_26  (
    .i0(inst_doa_i52_007),
    .i1(inst_doa_i53_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_26 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_27  (
    .i0(inst_doa_i54_007),
    .i1(inst_doa_i55_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_27 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_28  (
    .i0(inst_doa_i56_007),
    .i1(inst_doa_i57_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_28 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_29  (
    .i0(inst_doa_i58_007),
    .i1(inst_doa_i59_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_29 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_3  (
    .i0(inst_doa_i6_007),
    .i1(inst_doa_i7_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_3 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_30  (
    .i0(inst_doa_i60_007),
    .i1(inst_doa_i61_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_30 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_31  (
    .i0(inst_doa_i62_007),
    .i1(inst_doa_i63_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_31 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_4  (
    .i0(inst_doa_i8_007),
    .i1(inst_doa_i9_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_4 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_5  (
    .i0(inst_doa_i10_007),
    .i1(inst_doa_i11_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_5 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_6  (
    .i0(inst_doa_i12_007),
    .i1(inst_doa_i13_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_6 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_7  (
    .i0(inst_doa_i14_007),
    .i1(inst_doa_i15_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_7 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_8  (
    .i0(inst_doa_i16_007),
    .i1(inst_doa_i17_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_8 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_9  (
    .i0(inst_doa_i18_007),
    .i1(inst_doa_i19_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_9 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b7/B0_2 ),
    .i1(\inst_doa_mux_b7/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b7/B0_20 ),
    .i1(\inst_doa_mux_b7/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_10 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b7/B0_22 ),
    .i1(\inst_doa_mux_b7/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_11 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b7/B0_24 ),
    .i1(\inst_doa_mux_b7/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_12 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b7/B0_26 ),
    .i1(\inst_doa_mux_b7/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_13 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b7/B0_28 ),
    .i1(\inst_doa_mux_b7/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_14 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b7/B0_30 ),
    .i1(\inst_doa_mux_b7/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_15 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b7/B0_4 ),
    .i1(\inst_doa_mux_b7/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_2 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b7/B0_6 ),
    .i1(\inst_doa_mux_b7/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_3 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b7/B0_8 ),
    .i1(\inst_doa_mux_b7/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_4 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b7/B0_10 ),
    .i1(\inst_doa_mux_b7/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_5 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b7/B0_12 ),
    .i1(\inst_doa_mux_b7/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_6 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b7/B0_14 ),
    .i1(\inst_doa_mux_b7/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_7 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b7/B0_16 ),
    .i1(\inst_doa_mux_b7/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_8 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b7/B0_18 ),
    .i1(\inst_doa_mux_b7/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_9 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b7/B1_0 ),
    .i1(\inst_doa_mux_b7/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b7/B1_2 ),
    .i1(\inst_doa_mux_b7/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b7/B1_4 ),
    .i1(\inst_doa_mux_b7/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_2 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b7/B1_6 ),
    .i1(\inst_doa_mux_b7/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_3 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b7/B1_8 ),
    .i1(\inst_doa_mux_b7/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_4 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b7/B1_10 ),
    .i1(\inst_doa_mux_b7/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_5 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b7/B1_12 ),
    .i1(\inst_doa_mux_b7/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_6 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b7/B1_14 ),
    .i1(\inst_doa_mux_b7/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_7 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b7/B2_0 ),
    .i1(\inst_doa_mux_b7/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b7/B3_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b7/B2_2 ),
    .i1(\inst_doa_mux_b7/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b7/B3_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b7/B2_4 ),
    .i1(\inst_doa_mux_b7/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b7/B3_2 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b7/B2_6 ),
    .i1(\inst_doa_mux_b7/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b7/B3_3 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b7/B3_0 ),
    .i1(\inst_doa_mux_b7/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b7/B4_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b7/B3_2 ),
    .i1(\inst_doa_mux_b7/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b7/B4_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b7/B4_0 ),
    .i1(\inst_doa_mux_b7/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[7]));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_0  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i1_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_1  (
    .i0(inst_doa_i2_008),
    .i1(inst_doa_i3_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_10  (
    .i0(inst_doa_i20_008),
    .i1(inst_doa_i21_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_10 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_11  (
    .i0(inst_doa_i22_008),
    .i1(inst_doa_i23_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_11 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_12  (
    .i0(inst_doa_i24_008),
    .i1(inst_doa_i25_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_12 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_13  (
    .i0(inst_doa_i26_008),
    .i1(inst_doa_i27_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_13 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_14  (
    .i0(inst_doa_i28_008),
    .i1(inst_doa_i29_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_14 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_15  (
    .i0(inst_doa_i30_008),
    .i1(inst_doa_i31_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_15 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_16  (
    .i0(inst_doa_i32_008),
    .i1(inst_doa_i33_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_16 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_17  (
    .i0(inst_doa_i34_008),
    .i1(inst_doa_i35_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_17 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_18  (
    .i0(inst_doa_i36_008),
    .i1(inst_doa_i37_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_18 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_19  (
    .i0(inst_doa_i38_008),
    .i1(inst_doa_i39_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_19 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_2  (
    .i0(inst_doa_i4_008),
    .i1(inst_doa_i5_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_2 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_20  (
    .i0(inst_doa_i40_008),
    .i1(inst_doa_i41_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_20 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_21  (
    .i0(inst_doa_i42_008),
    .i1(inst_doa_i43_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_21 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_22  (
    .i0(inst_doa_i44_008),
    .i1(inst_doa_i45_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_22 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_23  (
    .i0(inst_doa_i46_008),
    .i1(inst_doa_i47_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_23 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_24  (
    .i0(inst_doa_i48_008),
    .i1(inst_doa_i49_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_24 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_25  (
    .i0(inst_doa_i50_008),
    .i1(inst_doa_i51_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_25 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_26  (
    .i0(inst_doa_i52_008),
    .i1(inst_doa_i53_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_26 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_27  (
    .i0(inst_doa_i54_008),
    .i1(inst_doa_i55_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_27 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_28  (
    .i0(inst_doa_i56_008),
    .i1(inst_doa_i57_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_28 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_29  (
    .i0(inst_doa_i58_008),
    .i1(inst_doa_i59_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_29 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_3  (
    .i0(inst_doa_i6_008),
    .i1(inst_doa_i7_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_3 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_30  (
    .i0(inst_doa_i60_008),
    .i1(inst_doa_i61_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_30 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_31  (
    .i0(inst_doa_i62_008),
    .i1(inst_doa_i63_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_31 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_4  (
    .i0(inst_doa_i8_008),
    .i1(inst_doa_i9_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_4 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_5  (
    .i0(inst_doa_i10_008),
    .i1(inst_doa_i11_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_5 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_6  (
    .i0(inst_doa_i12_008),
    .i1(inst_doa_i13_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_6 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_7  (
    .i0(inst_doa_i14_008),
    .i1(inst_doa_i15_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_7 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_8  (
    .i0(inst_doa_i16_008),
    .i1(inst_doa_i17_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_8 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_9  (
    .i0(inst_doa_i18_008),
    .i1(inst_doa_i19_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_9 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b8/B0_0 ),
    .i1(\inst_doa_mux_b8/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b8/B0_2 ),
    .i1(\inst_doa_mux_b8/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b8/B0_20 ),
    .i1(\inst_doa_mux_b8/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_10 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b8/B0_22 ),
    .i1(\inst_doa_mux_b8/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_11 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b8/B0_24 ),
    .i1(\inst_doa_mux_b8/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_12 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b8/B0_26 ),
    .i1(\inst_doa_mux_b8/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_13 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b8/B0_28 ),
    .i1(\inst_doa_mux_b8/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_14 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b8/B0_30 ),
    .i1(\inst_doa_mux_b8/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_15 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b8/B0_4 ),
    .i1(\inst_doa_mux_b8/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_2 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b8/B0_6 ),
    .i1(\inst_doa_mux_b8/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_3 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b8/B0_8 ),
    .i1(\inst_doa_mux_b8/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_4 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b8/B0_10 ),
    .i1(\inst_doa_mux_b8/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_5 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b8/B0_12 ),
    .i1(\inst_doa_mux_b8/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_6 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b8/B0_14 ),
    .i1(\inst_doa_mux_b8/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_7 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b8/B0_16 ),
    .i1(\inst_doa_mux_b8/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_8 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b8/B0_18 ),
    .i1(\inst_doa_mux_b8/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_9 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b8/B1_0 ),
    .i1(\inst_doa_mux_b8/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b8/B1_2 ),
    .i1(\inst_doa_mux_b8/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b8/B1_4 ),
    .i1(\inst_doa_mux_b8/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_2 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b8/B1_6 ),
    .i1(\inst_doa_mux_b8/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_3 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b8/B1_8 ),
    .i1(\inst_doa_mux_b8/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_4 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b8/B1_10 ),
    .i1(\inst_doa_mux_b8/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_5 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b8/B1_12 ),
    .i1(\inst_doa_mux_b8/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_6 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b8/B1_14 ),
    .i1(\inst_doa_mux_b8/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_7 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b8/B2_0 ),
    .i1(\inst_doa_mux_b8/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b8/B3_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b8/B2_2 ),
    .i1(\inst_doa_mux_b8/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b8/B3_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b8/B2_4 ),
    .i1(\inst_doa_mux_b8/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b8/B3_2 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b8/B2_6 ),
    .i1(\inst_doa_mux_b8/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b8/B3_3 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b8/B3_0 ),
    .i1(\inst_doa_mux_b8/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b8/B4_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b8/B3_2 ),
    .i1(\inst_doa_mux_b8/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b8/B4_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b8/B4_0 ),
    .i1(\inst_doa_mux_b8/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[8]));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

