module top( );



endmodule
