module Imgdata_send(
      input wire clk,
      input wire tft_de,
      input wire hcount,
      input wire vcount,
      output wire img_ack
  );
     

     
 endmodule