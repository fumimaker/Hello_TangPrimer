// Verilog netlist created by TD v4.2.217
// Sat Jul 28 11:33:58 2018

`timescale 1ns / 1ps
module img_cache  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_ram.v(14)
  (
  addra,
  addrb,
  cea,
  ceb,
  clka,
  clkb,
  dia,
  rsta,
  rstb,
  dob
  );

  input [15:0] addra;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_ram.v(23)
  input [15:0] addrb;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_ram.v(24)
  input cea;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_ram.v(25)
  input ceb;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_ram.v(26)
  input clka;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_ram.v(27)
  input clkb;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_ram.v(28)
  input [15:0] dia;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_ram.v(22)
  input rsta;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_ram.v(29)
  input rstb;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_ram.v(30)
  output [15:0] dob;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_ram.v(19)

  wire [0:6] addrb_piped;
  wire  \inst_dob_mux_b0/B0_0 ;
  wire  \inst_dob_mux_b0/B0_1 ;
  wire  \inst_dob_mux_b0/B0_10 ;
  wire  \inst_dob_mux_b0/B0_11 ;
  wire  \inst_dob_mux_b0/B0_12 ;
  wire  \inst_dob_mux_b0/B0_13 ;
  wire  \inst_dob_mux_b0/B0_14 ;
  wire  \inst_dob_mux_b0/B0_15 ;
  wire  \inst_dob_mux_b0/B0_16 ;
  wire  \inst_dob_mux_b0/B0_17 ;
  wire  \inst_dob_mux_b0/B0_18 ;
  wire  \inst_dob_mux_b0/B0_19 ;
  wire  \inst_dob_mux_b0/B0_2 ;
  wire  \inst_dob_mux_b0/B0_20 ;
  wire  \inst_dob_mux_b0/B0_21 ;
  wire  \inst_dob_mux_b0/B0_22 ;
  wire  \inst_dob_mux_b0/B0_23 ;
  wire  \inst_dob_mux_b0/B0_24 ;
  wire  \inst_dob_mux_b0/B0_25 ;
  wire  \inst_dob_mux_b0/B0_26 ;
  wire  \inst_dob_mux_b0/B0_27 ;
  wire  \inst_dob_mux_b0/B0_28 ;
  wire  \inst_dob_mux_b0/B0_29 ;
  wire  \inst_dob_mux_b0/B0_3 ;
  wire  \inst_dob_mux_b0/B0_30 ;
  wire  \inst_dob_mux_b0/B0_31 ;
  wire  \inst_dob_mux_b0/B0_32 ;
  wire  \inst_dob_mux_b0/B0_33 ;
  wire  \inst_dob_mux_b0/B0_34 ;
  wire  \inst_dob_mux_b0/B0_35 ;
  wire  \inst_dob_mux_b0/B0_36 ;
  wire  \inst_dob_mux_b0/B0_37 ;
  wire  \inst_dob_mux_b0/B0_38 ;
  wire  \inst_dob_mux_b0/B0_39 ;
  wire  \inst_dob_mux_b0/B0_4 ;
  wire  \inst_dob_mux_b0/B0_40 ;
  wire  \inst_dob_mux_b0/B0_41 ;
  wire  \inst_dob_mux_b0/B0_42 ;
  wire  \inst_dob_mux_b0/B0_43 ;
  wire  \inst_dob_mux_b0/B0_44 ;
  wire  \inst_dob_mux_b0/B0_45 ;
  wire  \inst_dob_mux_b0/B0_46 ;
  wire  \inst_dob_mux_b0/B0_47 ;
  wire  \inst_dob_mux_b0/B0_48 ;
  wire  \inst_dob_mux_b0/B0_49 ;
  wire  \inst_dob_mux_b0/B0_5 ;
  wire  \inst_dob_mux_b0/B0_50 ;
  wire  \inst_dob_mux_b0/B0_51 ;
  wire  \inst_dob_mux_b0/B0_52 ;
  wire  \inst_dob_mux_b0/B0_53 ;
  wire  \inst_dob_mux_b0/B0_54 ;
  wire  \inst_dob_mux_b0/B0_55 ;
  wire  \inst_dob_mux_b0/B0_56 ;
  wire  \inst_dob_mux_b0/B0_57 ;
  wire  \inst_dob_mux_b0/B0_58 ;
  wire  \inst_dob_mux_b0/B0_59 ;
  wire  \inst_dob_mux_b0/B0_6 ;
  wire  \inst_dob_mux_b0/B0_60 ;
  wire  \inst_dob_mux_b0/B0_61 ;
  wire  \inst_dob_mux_b0/B0_62 ;
  wire  \inst_dob_mux_b0/B0_63 ;
  wire  \inst_dob_mux_b0/B0_7 ;
  wire  \inst_dob_mux_b0/B0_8 ;
  wire  \inst_dob_mux_b0/B0_9 ;
  wire  \inst_dob_mux_b0/B1_0 ;
  wire  \inst_dob_mux_b0/B1_1 ;
  wire  \inst_dob_mux_b0/B1_10 ;
  wire  \inst_dob_mux_b0/B1_11 ;
  wire  \inst_dob_mux_b0/B1_12 ;
  wire  \inst_dob_mux_b0/B1_13 ;
  wire  \inst_dob_mux_b0/B1_14 ;
  wire  \inst_dob_mux_b0/B1_15 ;
  wire  \inst_dob_mux_b0/B1_16 ;
  wire  \inst_dob_mux_b0/B1_17 ;
  wire  \inst_dob_mux_b0/B1_18 ;
  wire  \inst_dob_mux_b0/B1_19 ;
  wire  \inst_dob_mux_b0/B1_2 ;
  wire  \inst_dob_mux_b0/B1_20 ;
  wire  \inst_dob_mux_b0/B1_21 ;
  wire  \inst_dob_mux_b0/B1_22 ;
  wire  \inst_dob_mux_b0/B1_23 ;
  wire  \inst_dob_mux_b0/B1_24 ;
  wire  \inst_dob_mux_b0/B1_25 ;
  wire  \inst_dob_mux_b0/B1_26 ;
  wire  \inst_dob_mux_b0/B1_27 ;
  wire  \inst_dob_mux_b0/B1_28 ;
  wire  \inst_dob_mux_b0/B1_29 ;
  wire  \inst_dob_mux_b0/B1_3 ;
  wire  \inst_dob_mux_b0/B1_30 ;
  wire  \inst_dob_mux_b0/B1_31 ;
  wire  \inst_dob_mux_b0/B1_4 ;
  wire  \inst_dob_mux_b0/B1_5 ;
  wire  \inst_dob_mux_b0/B1_6 ;
  wire  \inst_dob_mux_b0/B1_7 ;
  wire  \inst_dob_mux_b0/B1_8 ;
  wire  \inst_dob_mux_b0/B1_9 ;
  wire  \inst_dob_mux_b0/B2_0 ;
  wire  \inst_dob_mux_b0/B2_1 ;
  wire  \inst_dob_mux_b0/B2_10 ;
  wire  \inst_dob_mux_b0/B2_11 ;
  wire  \inst_dob_mux_b0/B2_12 ;
  wire  \inst_dob_mux_b0/B2_13 ;
  wire  \inst_dob_mux_b0/B2_14 ;
  wire  \inst_dob_mux_b0/B2_15 ;
  wire  \inst_dob_mux_b0/B2_2 ;
  wire  \inst_dob_mux_b0/B2_3 ;
  wire  \inst_dob_mux_b0/B2_4 ;
  wire  \inst_dob_mux_b0/B2_5 ;
  wire  \inst_dob_mux_b0/B2_6 ;
  wire  \inst_dob_mux_b0/B2_7 ;
  wire  \inst_dob_mux_b0/B2_8 ;
  wire  \inst_dob_mux_b0/B2_9 ;
  wire  \inst_dob_mux_b0/B3_0 ;
  wire  \inst_dob_mux_b0/B3_1 ;
  wire  \inst_dob_mux_b0/B3_2 ;
  wire  \inst_dob_mux_b0/B3_3 ;
  wire  \inst_dob_mux_b0/B3_4 ;
  wire  \inst_dob_mux_b0/B3_5 ;
  wire  \inst_dob_mux_b0/B3_6 ;
  wire  \inst_dob_mux_b0/B3_7 ;
  wire  \inst_dob_mux_b0/B4_0 ;
  wire  \inst_dob_mux_b0/B4_1 ;
  wire  \inst_dob_mux_b0/B4_2 ;
  wire  \inst_dob_mux_b0/B4_3 ;
  wire  \inst_dob_mux_b0/B5_0 ;
  wire  \inst_dob_mux_b0/B5_1 ;
  wire  \inst_dob_mux_b1/B0_0 ;
  wire  \inst_dob_mux_b1/B0_1 ;
  wire  \inst_dob_mux_b1/B0_10 ;
  wire  \inst_dob_mux_b1/B0_11 ;
  wire  \inst_dob_mux_b1/B0_12 ;
  wire  \inst_dob_mux_b1/B0_13 ;
  wire  \inst_dob_mux_b1/B0_14 ;
  wire  \inst_dob_mux_b1/B0_15 ;
  wire  \inst_dob_mux_b1/B0_16 ;
  wire  \inst_dob_mux_b1/B0_17 ;
  wire  \inst_dob_mux_b1/B0_18 ;
  wire  \inst_dob_mux_b1/B0_19 ;
  wire  \inst_dob_mux_b1/B0_2 ;
  wire  \inst_dob_mux_b1/B0_20 ;
  wire  \inst_dob_mux_b1/B0_21 ;
  wire  \inst_dob_mux_b1/B0_22 ;
  wire  \inst_dob_mux_b1/B0_23 ;
  wire  \inst_dob_mux_b1/B0_24 ;
  wire  \inst_dob_mux_b1/B0_25 ;
  wire  \inst_dob_mux_b1/B0_26 ;
  wire  \inst_dob_mux_b1/B0_27 ;
  wire  \inst_dob_mux_b1/B0_28 ;
  wire  \inst_dob_mux_b1/B0_29 ;
  wire  \inst_dob_mux_b1/B0_3 ;
  wire  \inst_dob_mux_b1/B0_30 ;
  wire  \inst_dob_mux_b1/B0_31 ;
  wire  \inst_dob_mux_b1/B0_32 ;
  wire  \inst_dob_mux_b1/B0_33 ;
  wire  \inst_dob_mux_b1/B0_34 ;
  wire  \inst_dob_mux_b1/B0_35 ;
  wire  \inst_dob_mux_b1/B0_36 ;
  wire  \inst_dob_mux_b1/B0_37 ;
  wire  \inst_dob_mux_b1/B0_38 ;
  wire  \inst_dob_mux_b1/B0_39 ;
  wire  \inst_dob_mux_b1/B0_4 ;
  wire  \inst_dob_mux_b1/B0_40 ;
  wire  \inst_dob_mux_b1/B0_41 ;
  wire  \inst_dob_mux_b1/B0_42 ;
  wire  \inst_dob_mux_b1/B0_43 ;
  wire  \inst_dob_mux_b1/B0_44 ;
  wire  \inst_dob_mux_b1/B0_45 ;
  wire  \inst_dob_mux_b1/B0_46 ;
  wire  \inst_dob_mux_b1/B0_47 ;
  wire  \inst_dob_mux_b1/B0_48 ;
  wire  \inst_dob_mux_b1/B0_49 ;
  wire  \inst_dob_mux_b1/B0_5 ;
  wire  \inst_dob_mux_b1/B0_50 ;
  wire  \inst_dob_mux_b1/B0_51 ;
  wire  \inst_dob_mux_b1/B0_52 ;
  wire  \inst_dob_mux_b1/B0_53 ;
  wire  \inst_dob_mux_b1/B0_54 ;
  wire  \inst_dob_mux_b1/B0_55 ;
  wire  \inst_dob_mux_b1/B0_56 ;
  wire  \inst_dob_mux_b1/B0_57 ;
  wire  \inst_dob_mux_b1/B0_58 ;
  wire  \inst_dob_mux_b1/B0_59 ;
  wire  \inst_dob_mux_b1/B0_6 ;
  wire  \inst_dob_mux_b1/B0_60 ;
  wire  \inst_dob_mux_b1/B0_61 ;
  wire  \inst_dob_mux_b1/B0_62 ;
  wire  \inst_dob_mux_b1/B0_63 ;
  wire  \inst_dob_mux_b1/B0_7 ;
  wire  \inst_dob_mux_b1/B0_8 ;
  wire  \inst_dob_mux_b1/B0_9 ;
  wire  \inst_dob_mux_b1/B1_0 ;
  wire  \inst_dob_mux_b1/B1_1 ;
  wire  \inst_dob_mux_b1/B1_10 ;
  wire  \inst_dob_mux_b1/B1_11 ;
  wire  \inst_dob_mux_b1/B1_12 ;
  wire  \inst_dob_mux_b1/B1_13 ;
  wire  \inst_dob_mux_b1/B1_14 ;
  wire  \inst_dob_mux_b1/B1_15 ;
  wire  \inst_dob_mux_b1/B1_16 ;
  wire  \inst_dob_mux_b1/B1_17 ;
  wire  \inst_dob_mux_b1/B1_18 ;
  wire  \inst_dob_mux_b1/B1_19 ;
  wire  \inst_dob_mux_b1/B1_2 ;
  wire  \inst_dob_mux_b1/B1_20 ;
  wire  \inst_dob_mux_b1/B1_21 ;
  wire  \inst_dob_mux_b1/B1_22 ;
  wire  \inst_dob_mux_b1/B1_23 ;
  wire  \inst_dob_mux_b1/B1_24 ;
  wire  \inst_dob_mux_b1/B1_25 ;
  wire  \inst_dob_mux_b1/B1_26 ;
  wire  \inst_dob_mux_b1/B1_27 ;
  wire  \inst_dob_mux_b1/B1_28 ;
  wire  \inst_dob_mux_b1/B1_29 ;
  wire  \inst_dob_mux_b1/B1_3 ;
  wire  \inst_dob_mux_b1/B1_30 ;
  wire  \inst_dob_mux_b1/B1_31 ;
  wire  \inst_dob_mux_b1/B1_4 ;
  wire  \inst_dob_mux_b1/B1_5 ;
  wire  \inst_dob_mux_b1/B1_6 ;
  wire  \inst_dob_mux_b1/B1_7 ;
  wire  \inst_dob_mux_b1/B1_8 ;
  wire  \inst_dob_mux_b1/B1_9 ;
  wire  \inst_dob_mux_b1/B2_0 ;
  wire  \inst_dob_mux_b1/B2_1 ;
  wire  \inst_dob_mux_b1/B2_10 ;
  wire  \inst_dob_mux_b1/B2_11 ;
  wire  \inst_dob_mux_b1/B2_12 ;
  wire  \inst_dob_mux_b1/B2_13 ;
  wire  \inst_dob_mux_b1/B2_14 ;
  wire  \inst_dob_mux_b1/B2_15 ;
  wire  \inst_dob_mux_b1/B2_2 ;
  wire  \inst_dob_mux_b1/B2_3 ;
  wire  \inst_dob_mux_b1/B2_4 ;
  wire  \inst_dob_mux_b1/B2_5 ;
  wire  \inst_dob_mux_b1/B2_6 ;
  wire  \inst_dob_mux_b1/B2_7 ;
  wire  \inst_dob_mux_b1/B2_8 ;
  wire  \inst_dob_mux_b1/B2_9 ;
  wire  \inst_dob_mux_b1/B3_0 ;
  wire  \inst_dob_mux_b1/B3_1 ;
  wire  \inst_dob_mux_b1/B3_2 ;
  wire  \inst_dob_mux_b1/B3_3 ;
  wire  \inst_dob_mux_b1/B3_4 ;
  wire  \inst_dob_mux_b1/B3_5 ;
  wire  \inst_dob_mux_b1/B3_6 ;
  wire  \inst_dob_mux_b1/B3_7 ;
  wire  \inst_dob_mux_b1/B4_0 ;
  wire  \inst_dob_mux_b1/B4_1 ;
  wire  \inst_dob_mux_b1/B4_2 ;
  wire  \inst_dob_mux_b1/B4_3 ;
  wire  \inst_dob_mux_b1/B5_0 ;
  wire  \inst_dob_mux_b1/B5_1 ;
  wire  \inst_dob_mux_b10/B0_0 ;
  wire  \inst_dob_mux_b10/B0_1 ;
  wire  \inst_dob_mux_b10/B0_10 ;
  wire  \inst_dob_mux_b10/B0_11 ;
  wire  \inst_dob_mux_b10/B0_12 ;
  wire  \inst_dob_mux_b10/B0_13 ;
  wire  \inst_dob_mux_b10/B0_14 ;
  wire  \inst_dob_mux_b10/B0_15 ;
  wire  \inst_dob_mux_b10/B0_16 ;
  wire  \inst_dob_mux_b10/B0_17 ;
  wire  \inst_dob_mux_b10/B0_18 ;
  wire  \inst_dob_mux_b10/B0_19 ;
  wire  \inst_dob_mux_b10/B0_2 ;
  wire  \inst_dob_mux_b10/B0_20 ;
  wire  \inst_dob_mux_b10/B0_21 ;
  wire  \inst_dob_mux_b10/B0_22 ;
  wire  \inst_dob_mux_b10/B0_23 ;
  wire  \inst_dob_mux_b10/B0_24 ;
  wire  \inst_dob_mux_b10/B0_25 ;
  wire  \inst_dob_mux_b10/B0_26 ;
  wire  \inst_dob_mux_b10/B0_27 ;
  wire  \inst_dob_mux_b10/B0_28 ;
  wire  \inst_dob_mux_b10/B0_29 ;
  wire  \inst_dob_mux_b10/B0_3 ;
  wire  \inst_dob_mux_b10/B0_30 ;
  wire  \inst_dob_mux_b10/B0_31 ;
  wire  \inst_dob_mux_b10/B0_32 ;
  wire  \inst_dob_mux_b10/B0_33 ;
  wire  \inst_dob_mux_b10/B0_34 ;
  wire  \inst_dob_mux_b10/B0_35 ;
  wire  \inst_dob_mux_b10/B0_36 ;
  wire  \inst_dob_mux_b10/B0_37 ;
  wire  \inst_dob_mux_b10/B0_38 ;
  wire  \inst_dob_mux_b10/B0_39 ;
  wire  \inst_dob_mux_b10/B0_4 ;
  wire  \inst_dob_mux_b10/B0_40 ;
  wire  \inst_dob_mux_b10/B0_41 ;
  wire  \inst_dob_mux_b10/B0_42 ;
  wire  \inst_dob_mux_b10/B0_43 ;
  wire  \inst_dob_mux_b10/B0_44 ;
  wire  \inst_dob_mux_b10/B0_45 ;
  wire  \inst_dob_mux_b10/B0_46 ;
  wire  \inst_dob_mux_b10/B0_47 ;
  wire  \inst_dob_mux_b10/B0_48 ;
  wire  \inst_dob_mux_b10/B0_49 ;
  wire  \inst_dob_mux_b10/B0_5 ;
  wire  \inst_dob_mux_b10/B0_50 ;
  wire  \inst_dob_mux_b10/B0_51 ;
  wire  \inst_dob_mux_b10/B0_52 ;
  wire  \inst_dob_mux_b10/B0_53 ;
  wire  \inst_dob_mux_b10/B0_54 ;
  wire  \inst_dob_mux_b10/B0_55 ;
  wire  \inst_dob_mux_b10/B0_56 ;
  wire  \inst_dob_mux_b10/B0_57 ;
  wire  \inst_dob_mux_b10/B0_58 ;
  wire  \inst_dob_mux_b10/B0_59 ;
  wire  \inst_dob_mux_b10/B0_6 ;
  wire  \inst_dob_mux_b10/B0_60 ;
  wire  \inst_dob_mux_b10/B0_61 ;
  wire  \inst_dob_mux_b10/B0_62 ;
  wire  \inst_dob_mux_b10/B0_63 ;
  wire  \inst_dob_mux_b10/B0_7 ;
  wire  \inst_dob_mux_b10/B0_8 ;
  wire  \inst_dob_mux_b10/B0_9 ;
  wire  \inst_dob_mux_b10/B1_0 ;
  wire  \inst_dob_mux_b10/B1_1 ;
  wire  \inst_dob_mux_b10/B1_10 ;
  wire  \inst_dob_mux_b10/B1_11 ;
  wire  \inst_dob_mux_b10/B1_12 ;
  wire  \inst_dob_mux_b10/B1_13 ;
  wire  \inst_dob_mux_b10/B1_14 ;
  wire  \inst_dob_mux_b10/B1_15 ;
  wire  \inst_dob_mux_b10/B1_16 ;
  wire  \inst_dob_mux_b10/B1_17 ;
  wire  \inst_dob_mux_b10/B1_18 ;
  wire  \inst_dob_mux_b10/B1_19 ;
  wire  \inst_dob_mux_b10/B1_2 ;
  wire  \inst_dob_mux_b10/B1_20 ;
  wire  \inst_dob_mux_b10/B1_21 ;
  wire  \inst_dob_mux_b10/B1_22 ;
  wire  \inst_dob_mux_b10/B1_23 ;
  wire  \inst_dob_mux_b10/B1_24 ;
  wire  \inst_dob_mux_b10/B1_25 ;
  wire  \inst_dob_mux_b10/B1_26 ;
  wire  \inst_dob_mux_b10/B1_27 ;
  wire  \inst_dob_mux_b10/B1_28 ;
  wire  \inst_dob_mux_b10/B1_29 ;
  wire  \inst_dob_mux_b10/B1_3 ;
  wire  \inst_dob_mux_b10/B1_30 ;
  wire  \inst_dob_mux_b10/B1_31 ;
  wire  \inst_dob_mux_b10/B1_4 ;
  wire  \inst_dob_mux_b10/B1_5 ;
  wire  \inst_dob_mux_b10/B1_6 ;
  wire  \inst_dob_mux_b10/B1_7 ;
  wire  \inst_dob_mux_b10/B1_8 ;
  wire  \inst_dob_mux_b10/B1_9 ;
  wire  \inst_dob_mux_b10/B2_0 ;
  wire  \inst_dob_mux_b10/B2_1 ;
  wire  \inst_dob_mux_b10/B2_10 ;
  wire  \inst_dob_mux_b10/B2_11 ;
  wire  \inst_dob_mux_b10/B2_12 ;
  wire  \inst_dob_mux_b10/B2_13 ;
  wire  \inst_dob_mux_b10/B2_14 ;
  wire  \inst_dob_mux_b10/B2_15 ;
  wire  \inst_dob_mux_b10/B2_2 ;
  wire  \inst_dob_mux_b10/B2_3 ;
  wire  \inst_dob_mux_b10/B2_4 ;
  wire  \inst_dob_mux_b10/B2_5 ;
  wire  \inst_dob_mux_b10/B2_6 ;
  wire  \inst_dob_mux_b10/B2_7 ;
  wire  \inst_dob_mux_b10/B2_8 ;
  wire  \inst_dob_mux_b10/B2_9 ;
  wire  \inst_dob_mux_b10/B3_0 ;
  wire  \inst_dob_mux_b10/B3_1 ;
  wire  \inst_dob_mux_b10/B3_2 ;
  wire  \inst_dob_mux_b10/B3_3 ;
  wire  \inst_dob_mux_b10/B3_4 ;
  wire  \inst_dob_mux_b10/B3_5 ;
  wire  \inst_dob_mux_b10/B3_6 ;
  wire  \inst_dob_mux_b10/B3_7 ;
  wire  \inst_dob_mux_b10/B4_0 ;
  wire  \inst_dob_mux_b10/B4_1 ;
  wire  \inst_dob_mux_b10/B4_2 ;
  wire  \inst_dob_mux_b10/B4_3 ;
  wire  \inst_dob_mux_b10/B5_0 ;
  wire  \inst_dob_mux_b10/B5_1 ;
  wire  \inst_dob_mux_b11/B0_0 ;
  wire  \inst_dob_mux_b11/B0_1 ;
  wire  \inst_dob_mux_b11/B0_10 ;
  wire  \inst_dob_mux_b11/B0_11 ;
  wire  \inst_dob_mux_b11/B0_12 ;
  wire  \inst_dob_mux_b11/B0_13 ;
  wire  \inst_dob_mux_b11/B0_14 ;
  wire  \inst_dob_mux_b11/B0_15 ;
  wire  \inst_dob_mux_b11/B0_16 ;
  wire  \inst_dob_mux_b11/B0_17 ;
  wire  \inst_dob_mux_b11/B0_18 ;
  wire  \inst_dob_mux_b11/B0_19 ;
  wire  \inst_dob_mux_b11/B0_2 ;
  wire  \inst_dob_mux_b11/B0_20 ;
  wire  \inst_dob_mux_b11/B0_21 ;
  wire  \inst_dob_mux_b11/B0_22 ;
  wire  \inst_dob_mux_b11/B0_23 ;
  wire  \inst_dob_mux_b11/B0_24 ;
  wire  \inst_dob_mux_b11/B0_25 ;
  wire  \inst_dob_mux_b11/B0_26 ;
  wire  \inst_dob_mux_b11/B0_27 ;
  wire  \inst_dob_mux_b11/B0_28 ;
  wire  \inst_dob_mux_b11/B0_29 ;
  wire  \inst_dob_mux_b11/B0_3 ;
  wire  \inst_dob_mux_b11/B0_30 ;
  wire  \inst_dob_mux_b11/B0_31 ;
  wire  \inst_dob_mux_b11/B0_32 ;
  wire  \inst_dob_mux_b11/B0_33 ;
  wire  \inst_dob_mux_b11/B0_34 ;
  wire  \inst_dob_mux_b11/B0_35 ;
  wire  \inst_dob_mux_b11/B0_36 ;
  wire  \inst_dob_mux_b11/B0_37 ;
  wire  \inst_dob_mux_b11/B0_38 ;
  wire  \inst_dob_mux_b11/B0_39 ;
  wire  \inst_dob_mux_b11/B0_4 ;
  wire  \inst_dob_mux_b11/B0_40 ;
  wire  \inst_dob_mux_b11/B0_41 ;
  wire  \inst_dob_mux_b11/B0_42 ;
  wire  \inst_dob_mux_b11/B0_43 ;
  wire  \inst_dob_mux_b11/B0_44 ;
  wire  \inst_dob_mux_b11/B0_45 ;
  wire  \inst_dob_mux_b11/B0_46 ;
  wire  \inst_dob_mux_b11/B0_47 ;
  wire  \inst_dob_mux_b11/B0_48 ;
  wire  \inst_dob_mux_b11/B0_49 ;
  wire  \inst_dob_mux_b11/B0_5 ;
  wire  \inst_dob_mux_b11/B0_50 ;
  wire  \inst_dob_mux_b11/B0_51 ;
  wire  \inst_dob_mux_b11/B0_52 ;
  wire  \inst_dob_mux_b11/B0_53 ;
  wire  \inst_dob_mux_b11/B0_54 ;
  wire  \inst_dob_mux_b11/B0_55 ;
  wire  \inst_dob_mux_b11/B0_56 ;
  wire  \inst_dob_mux_b11/B0_57 ;
  wire  \inst_dob_mux_b11/B0_58 ;
  wire  \inst_dob_mux_b11/B0_59 ;
  wire  \inst_dob_mux_b11/B0_6 ;
  wire  \inst_dob_mux_b11/B0_60 ;
  wire  \inst_dob_mux_b11/B0_61 ;
  wire  \inst_dob_mux_b11/B0_62 ;
  wire  \inst_dob_mux_b11/B0_63 ;
  wire  \inst_dob_mux_b11/B0_7 ;
  wire  \inst_dob_mux_b11/B0_8 ;
  wire  \inst_dob_mux_b11/B0_9 ;
  wire  \inst_dob_mux_b11/B1_0 ;
  wire  \inst_dob_mux_b11/B1_1 ;
  wire  \inst_dob_mux_b11/B1_10 ;
  wire  \inst_dob_mux_b11/B1_11 ;
  wire  \inst_dob_mux_b11/B1_12 ;
  wire  \inst_dob_mux_b11/B1_13 ;
  wire  \inst_dob_mux_b11/B1_14 ;
  wire  \inst_dob_mux_b11/B1_15 ;
  wire  \inst_dob_mux_b11/B1_16 ;
  wire  \inst_dob_mux_b11/B1_17 ;
  wire  \inst_dob_mux_b11/B1_18 ;
  wire  \inst_dob_mux_b11/B1_19 ;
  wire  \inst_dob_mux_b11/B1_2 ;
  wire  \inst_dob_mux_b11/B1_20 ;
  wire  \inst_dob_mux_b11/B1_21 ;
  wire  \inst_dob_mux_b11/B1_22 ;
  wire  \inst_dob_mux_b11/B1_23 ;
  wire  \inst_dob_mux_b11/B1_24 ;
  wire  \inst_dob_mux_b11/B1_25 ;
  wire  \inst_dob_mux_b11/B1_26 ;
  wire  \inst_dob_mux_b11/B1_27 ;
  wire  \inst_dob_mux_b11/B1_28 ;
  wire  \inst_dob_mux_b11/B1_29 ;
  wire  \inst_dob_mux_b11/B1_3 ;
  wire  \inst_dob_mux_b11/B1_30 ;
  wire  \inst_dob_mux_b11/B1_31 ;
  wire  \inst_dob_mux_b11/B1_4 ;
  wire  \inst_dob_mux_b11/B1_5 ;
  wire  \inst_dob_mux_b11/B1_6 ;
  wire  \inst_dob_mux_b11/B1_7 ;
  wire  \inst_dob_mux_b11/B1_8 ;
  wire  \inst_dob_mux_b11/B1_9 ;
  wire  \inst_dob_mux_b11/B2_0 ;
  wire  \inst_dob_mux_b11/B2_1 ;
  wire  \inst_dob_mux_b11/B2_10 ;
  wire  \inst_dob_mux_b11/B2_11 ;
  wire  \inst_dob_mux_b11/B2_12 ;
  wire  \inst_dob_mux_b11/B2_13 ;
  wire  \inst_dob_mux_b11/B2_14 ;
  wire  \inst_dob_mux_b11/B2_15 ;
  wire  \inst_dob_mux_b11/B2_2 ;
  wire  \inst_dob_mux_b11/B2_3 ;
  wire  \inst_dob_mux_b11/B2_4 ;
  wire  \inst_dob_mux_b11/B2_5 ;
  wire  \inst_dob_mux_b11/B2_6 ;
  wire  \inst_dob_mux_b11/B2_7 ;
  wire  \inst_dob_mux_b11/B2_8 ;
  wire  \inst_dob_mux_b11/B2_9 ;
  wire  \inst_dob_mux_b11/B3_0 ;
  wire  \inst_dob_mux_b11/B3_1 ;
  wire  \inst_dob_mux_b11/B3_2 ;
  wire  \inst_dob_mux_b11/B3_3 ;
  wire  \inst_dob_mux_b11/B3_4 ;
  wire  \inst_dob_mux_b11/B3_5 ;
  wire  \inst_dob_mux_b11/B3_6 ;
  wire  \inst_dob_mux_b11/B3_7 ;
  wire  \inst_dob_mux_b11/B4_0 ;
  wire  \inst_dob_mux_b11/B4_1 ;
  wire  \inst_dob_mux_b11/B4_2 ;
  wire  \inst_dob_mux_b11/B4_3 ;
  wire  \inst_dob_mux_b11/B5_0 ;
  wire  \inst_dob_mux_b11/B5_1 ;
  wire  \inst_dob_mux_b12/B0_0 ;
  wire  \inst_dob_mux_b12/B0_1 ;
  wire  \inst_dob_mux_b12/B0_10 ;
  wire  \inst_dob_mux_b12/B0_11 ;
  wire  \inst_dob_mux_b12/B0_12 ;
  wire  \inst_dob_mux_b12/B0_13 ;
  wire  \inst_dob_mux_b12/B0_14 ;
  wire  \inst_dob_mux_b12/B0_15 ;
  wire  \inst_dob_mux_b12/B0_16 ;
  wire  \inst_dob_mux_b12/B0_17 ;
  wire  \inst_dob_mux_b12/B0_18 ;
  wire  \inst_dob_mux_b12/B0_19 ;
  wire  \inst_dob_mux_b12/B0_2 ;
  wire  \inst_dob_mux_b12/B0_20 ;
  wire  \inst_dob_mux_b12/B0_21 ;
  wire  \inst_dob_mux_b12/B0_22 ;
  wire  \inst_dob_mux_b12/B0_23 ;
  wire  \inst_dob_mux_b12/B0_24 ;
  wire  \inst_dob_mux_b12/B0_25 ;
  wire  \inst_dob_mux_b12/B0_26 ;
  wire  \inst_dob_mux_b12/B0_27 ;
  wire  \inst_dob_mux_b12/B0_28 ;
  wire  \inst_dob_mux_b12/B0_29 ;
  wire  \inst_dob_mux_b12/B0_3 ;
  wire  \inst_dob_mux_b12/B0_30 ;
  wire  \inst_dob_mux_b12/B0_31 ;
  wire  \inst_dob_mux_b12/B0_32 ;
  wire  \inst_dob_mux_b12/B0_33 ;
  wire  \inst_dob_mux_b12/B0_34 ;
  wire  \inst_dob_mux_b12/B0_35 ;
  wire  \inst_dob_mux_b12/B0_36 ;
  wire  \inst_dob_mux_b12/B0_37 ;
  wire  \inst_dob_mux_b12/B0_38 ;
  wire  \inst_dob_mux_b12/B0_39 ;
  wire  \inst_dob_mux_b12/B0_4 ;
  wire  \inst_dob_mux_b12/B0_40 ;
  wire  \inst_dob_mux_b12/B0_41 ;
  wire  \inst_dob_mux_b12/B0_42 ;
  wire  \inst_dob_mux_b12/B0_43 ;
  wire  \inst_dob_mux_b12/B0_44 ;
  wire  \inst_dob_mux_b12/B0_45 ;
  wire  \inst_dob_mux_b12/B0_46 ;
  wire  \inst_dob_mux_b12/B0_47 ;
  wire  \inst_dob_mux_b12/B0_48 ;
  wire  \inst_dob_mux_b12/B0_49 ;
  wire  \inst_dob_mux_b12/B0_5 ;
  wire  \inst_dob_mux_b12/B0_50 ;
  wire  \inst_dob_mux_b12/B0_51 ;
  wire  \inst_dob_mux_b12/B0_52 ;
  wire  \inst_dob_mux_b12/B0_53 ;
  wire  \inst_dob_mux_b12/B0_54 ;
  wire  \inst_dob_mux_b12/B0_55 ;
  wire  \inst_dob_mux_b12/B0_56 ;
  wire  \inst_dob_mux_b12/B0_57 ;
  wire  \inst_dob_mux_b12/B0_58 ;
  wire  \inst_dob_mux_b12/B0_59 ;
  wire  \inst_dob_mux_b12/B0_6 ;
  wire  \inst_dob_mux_b12/B0_60 ;
  wire  \inst_dob_mux_b12/B0_61 ;
  wire  \inst_dob_mux_b12/B0_62 ;
  wire  \inst_dob_mux_b12/B0_63 ;
  wire  \inst_dob_mux_b12/B0_7 ;
  wire  \inst_dob_mux_b12/B0_8 ;
  wire  \inst_dob_mux_b12/B0_9 ;
  wire  \inst_dob_mux_b12/B1_0 ;
  wire  \inst_dob_mux_b12/B1_1 ;
  wire  \inst_dob_mux_b12/B1_10 ;
  wire  \inst_dob_mux_b12/B1_11 ;
  wire  \inst_dob_mux_b12/B1_12 ;
  wire  \inst_dob_mux_b12/B1_13 ;
  wire  \inst_dob_mux_b12/B1_14 ;
  wire  \inst_dob_mux_b12/B1_15 ;
  wire  \inst_dob_mux_b12/B1_16 ;
  wire  \inst_dob_mux_b12/B1_17 ;
  wire  \inst_dob_mux_b12/B1_18 ;
  wire  \inst_dob_mux_b12/B1_19 ;
  wire  \inst_dob_mux_b12/B1_2 ;
  wire  \inst_dob_mux_b12/B1_20 ;
  wire  \inst_dob_mux_b12/B1_21 ;
  wire  \inst_dob_mux_b12/B1_22 ;
  wire  \inst_dob_mux_b12/B1_23 ;
  wire  \inst_dob_mux_b12/B1_24 ;
  wire  \inst_dob_mux_b12/B1_25 ;
  wire  \inst_dob_mux_b12/B1_26 ;
  wire  \inst_dob_mux_b12/B1_27 ;
  wire  \inst_dob_mux_b12/B1_28 ;
  wire  \inst_dob_mux_b12/B1_29 ;
  wire  \inst_dob_mux_b12/B1_3 ;
  wire  \inst_dob_mux_b12/B1_30 ;
  wire  \inst_dob_mux_b12/B1_31 ;
  wire  \inst_dob_mux_b12/B1_4 ;
  wire  \inst_dob_mux_b12/B1_5 ;
  wire  \inst_dob_mux_b12/B1_6 ;
  wire  \inst_dob_mux_b12/B1_7 ;
  wire  \inst_dob_mux_b12/B1_8 ;
  wire  \inst_dob_mux_b12/B1_9 ;
  wire  \inst_dob_mux_b12/B2_0 ;
  wire  \inst_dob_mux_b12/B2_1 ;
  wire  \inst_dob_mux_b12/B2_10 ;
  wire  \inst_dob_mux_b12/B2_11 ;
  wire  \inst_dob_mux_b12/B2_12 ;
  wire  \inst_dob_mux_b12/B2_13 ;
  wire  \inst_dob_mux_b12/B2_14 ;
  wire  \inst_dob_mux_b12/B2_15 ;
  wire  \inst_dob_mux_b12/B2_2 ;
  wire  \inst_dob_mux_b12/B2_3 ;
  wire  \inst_dob_mux_b12/B2_4 ;
  wire  \inst_dob_mux_b12/B2_5 ;
  wire  \inst_dob_mux_b12/B2_6 ;
  wire  \inst_dob_mux_b12/B2_7 ;
  wire  \inst_dob_mux_b12/B2_8 ;
  wire  \inst_dob_mux_b12/B2_9 ;
  wire  \inst_dob_mux_b12/B3_0 ;
  wire  \inst_dob_mux_b12/B3_1 ;
  wire  \inst_dob_mux_b12/B3_2 ;
  wire  \inst_dob_mux_b12/B3_3 ;
  wire  \inst_dob_mux_b12/B3_4 ;
  wire  \inst_dob_mux_b12/B3_5 ;
  wire  \inst_dob_mux_b12/B3_6 ;
  wire  \inst_dob_mux_b12/B3_7 ;
  wire  \inst_dob_mux_b12/B4_0 ;
  wire  \inst_dob_mux_b12/B4_1 ;
  wire  \inst_dob_mux_b12/B4_2 ;
  wire  \inst_dob_mux_b12/B4_3 ;
  wire  \inst_dob_mux_b12/B5_0 ;
  wire  \inst_dob_mux_b12/B5_1 ;
  wire  \inst_dob_mux_b13/B0_0 ;
  wire  \inst_dob_mux_b13/B0_1 ;
  wire  \inst_dob_mux_b13/B0_10 ;
  wire  \inst_dob_mux_b13/B0_11 ;
  wire  \inst_dob_mux_b13/B0_12 ;
  wire  \inst_dob_mux_b13/B0_13 ;
  wire  \inst_dob_mux_b13/B0_14 ;
  wire  \inst_dob_mux_b13/B0_15 ;
  wire  \inst_dob_mux_b13/B0_16 ;
  wire  \inst_dob_mux_b13/B0_17 ;
  wire  \inst_dob_mux_b13/B0_18 ;
  wire  \inst_dob_mux_b13/B0_19 ;
  wire  \inst_dob_mux_b13/B0_2 ;
  wire  \inst_dob_mux_b13/B0_20 ;
  wire  \inst_dob_mux_b13/B0_21 ;
  wire  \inst_dob_mux_b13/B0_22 ;
  wire  \inst_dob_mux_b13/B0_23 ;
  wire  \inst_dob_mux_b13/B0_24 ;
  wire  \inst_dob_mux_b13/B0_25 ;
  wire  \inst_dob_mux_b13/B0_26 ;
  wire  \inst_dob_mux_b13/B0_27 ;
  wire  \inst_dob_mux_b13/B0_28 ;
  wire  \inst_dob_mux_b13/B0_29 ;
  wire  \inst_dob_mux_b13/B0_3 ;
  wire  \inst_dob_mux_b13/B0_30 ;
  wire  \inst_dob_mux_b13/B0_31 ;
  wire  \inst_dob_mux_b13/B0_32 ;
  wire  \inst_dob_mux_b13/B0_33 ;
  wire  \inst_dob_mux_b13/B0_34 ;
  wire  \inst_dob_mux_b13/B0_35 ;
  wire  \inst_dob_mux_b13/B0_36 ;
  wire  \inst_dob_mux_b13/B0_37 ;
  wire  \inst_dob_mux_b13/B0_38 ;
  wire  \inst_dob_mux_b13/B0_39 ;
  wire  \inst_dob_mux_b13/B0_4 ;
  wire  \inst_dob_mux_b13/B0_40 ;
  wire  \inst_dob_mux_b13/B0_41 ;
  wire  \inst_dob_mux_b13/B0_42 ;
  wire  \inst_dob_mux_b13/B0_43 ;
  wire  \inst_dob_mux_b13/B0_44 ;
  wire  \inst_dob_mux_b13/B0_45 ;
  wire  \inst_dob_mux_b13/B0_46 ;
  wire  \inst_dob_mux_b13/B0_47 ;
  wire  \inst_dob_mux_b13/B0_48 ;
  wire  \inst_dob_mux_b13/B0_49 ;
  wire  \inst_dob_mux_b13/B0_5 ;
  wire  \inst_dob_mux_b13/B0_50 ;
  wire  \inst_dob_mux_b13/B0_51 ;
  wire  \inst_dob_mux_b13/B0_52 ;
  wire  \inst_dob_mux_b13/B0_53 ;
  wire  \inst_dob_mux_b13/B0_54 ;
  wire  \inst_dob_mux_b13/B0_55 ;
  wire  \inst_dob_mux_b13/B0_56 ;
  wire  \inst_dob_mux_b13/B0_57 ;
  wire  \inst_dob_mux_b13/B0_58 ;
  wire  \inst_dob_mux_b13/B0_59 ;
  wire  \inst_dob_mux_b13/B0_6 ;
  wire  \inst_dob_mux_b13/B0_60 ;
  wire  \inst_dob_mux_b13/B0_61 ;
  wire  \inst_dob_mux_b13/B0_62 ;
  wire  \inst_dob_mux_b13/B0_63 ;
  wire  \inst_dob_mux_b13/B0_7 ;
  wire  \inst_dob_mux_b13/B0_8 ;
  wire  \inst_dob_mux_b13/B0_9 ;
  wire  \inst_dob_mux_b13/B1_0 ;
  wire  \inst_dob_mux_b13/B1_1 ;
  wire  \inst_dob_mux_b13/B1_10 ;
  wire  \inst_dob_mux_b13/B1_11 ;
  wire  \inst_dob_mux_b13/B1_12 ;
  wire  \inst_dob_mux_b13/B1_13 ;
  wire  \inst_dob_mux_b13/B1_14 ;
  wire  \inst_dob_mux_b13/B1_15 ;
  wire  \inst_dob_mux_b13/B1_16 ;
  wire  \inst_dob_mux_b13/B1_17 ;
  wire  \inst_dob_mux_b13/B1_18 ;
  wire  \inst_dob_mux_b13/B1_19 ;
  wire  \inst_dob_mux_b13/B1_2 ;
  wire  \inst_dob_mux_b13/B1_20 ;
  wire  \inst_dob_mux_b13/B1_21 ;
  wire  \inst_dob_mux_b13/B1_22 ;
  wire  \inst_dob_mux_b13/B1_23 ;
  wire  \inst_dob_mux_b13/B1_24 ;
  wire  \inst_dob_mux_b13/B1_25 ;
  wire  \inst_dob_mux_b13/B1_26 ;
  wire  \inst_dob_mux_b13/B1_27 ;
  wire  \inst_dob_mux_b13/B1_28 ;
  wire  \inst_dob_mux_b13/B1_29 ;
  wire  \inst_dob_mux_b13/B1_3 ;
  wire  \inst_dob_mux_b13/B1_30 ;
  wire  \inst_dob_mux_b13/B1_31 ;
  wire  \inst_dob_mux_b13/B1_4 ;
  wire  \inst_dob_mux_b13/B1_5 ;
  wire  \inst_dob_mux_b13/B1_6 ;
  wire  \inst_dob_mux_b13/B1_7 ;
  wire  \inst_dob_mux_b13/B1_8 ;
  wire  \inst_dob_mux_b13/B1_9 ;
  wire  \inst_dob_mux_b13/B2_0 ;
  wire  \inst_dob_mux_b13/B2_1 ;
  wire  \inst_dob_mux_b13/B2_10 ;
  wire  \inst_dob_mux_b13/B2_11 ;
  wire  \inst_dob_mux_b13/B2_12 ;
  wire  \inst_dob_mux_b13/B2_13 ;
  wire  \inst_dob_mux_b13/B2_14 ;
  wire  \inst_dob_mux_b13/B2_15 ;
  wire  \inst_dob_mux_b13/B2_2 ;
  wire  \inst_dob_mux_b13/B2_3 ;
  wire  \inst_dob_mux_b13/B2_4 ;
  wire  \inst_dob_mux_b13/B2_5 ;
  wire  \inst_dob_mux_b13/B2_6 ;
  wire  \inst_dob_mux_b13/B2_7 ;
  wire  \inst_dob_mux_b13/B2_8 ;
  wire  \inst_dob_mux_b13/B2_9 ;
  wire  \inst_dob_mux_b13/B3_0 ;
  wire  \inst_dob_mux_b13/B3_1 ;
  wire  \inst_dob_mux_b13/B3_2 ;
  wire  \inst_dob_mux_b13/B3_3 ;
  wire  \inst_dob_mux_b13/B3_4 ;
  wire  \inst_dob_mux_b13/B3_5 ;
  wire  \inst_dob_mux_b13/B3_6 ;
  wire  \inst_dob_mux_b13/B3_7 ;
  wire  \inst_dob_mux_b13/B4_0 ;
  wire  \inst_dob_mux_b13/B4_1 ;
  wire  \inst_dob_mux_b13/B4_2 ;
  wire  \inst_dob_mux_b13/B4_3 ;
  wire  \inst_dob_mux_b13/B5_0 ;
  wire  \inst_dob_mux_b13/B5_1 ;
  wire  \inst_dob_mux_b14/B0_0 ;
  wire  \inst_dob_mux_b14/B0_1 ;
  wire  \inst_dob_mux_b14/B0_10 ;
  wire  \inst_dob_mux_b14/B0_11 ;
  wire  \inst_dob_mux_b14/B0_12 ;
  wire  \inst_dob_mux_b14/B0_13 ;
  wire  \inst_dob_mux_b14/B0_14 ;
  wire  \inst_dob_mux_b14/B0_15 ;
  wire  \inst_dob_mux_b14/B0_16 ;
  wire  \inst_dob_mux_b14/B0_17 ;
  wire  \inst_dob_mux_b14/B0_18 ;
  wire  \inst_dob_mux_b14/B0_19 ;
  wire  \inst_dob_mux_b14/B0_2 ;
  wire  \inst_dob_mux_b14/B0_20 ;
  wire  \inst_dob_mux_b14/B0_21 ;
  wire  \inst_dob_mux_b14/B0_22 ;
  wire  \inst_dob_mux_b14/B0_23 ;
  wire  \inst_dob_mux_b14/B0_24 ;
  wire  \inst_dob_mux_b14/B0_25 ;
  wire  \inst_dob_mux_b14/B0_26 ;
  wire  \inst_dob_mux_b14/B0_27 ;
  wire  \inst_dob_mux_b14/B0_28 ;
  wire  \inst_dob_mux_b14/B0_29 ;
  wire  \inst_dob_mux_b14/B0_3 ;
  wire  \inst_dob_mux_b14/B0_30 ;
  wire  \inst_dob_mux_b14/B0_31 ;
  wire  \inst_dob_mux_b14/B0_32 ;
  wire  \inst_dob_mux_b14/B0_33 ;
  wire  \inst_dob_mux_b14/B0_34 ;
  wire  \inst_dob_mux_b14/B0_35 ;
  wire  \inst_dob_mux_b14/B0_36 ;
  wire  \inst_dob_mux_b14/B0_37 ;
  wire  \inst_dob_mux_b14/B0_38 ;
  wire  \inst_dob_mux_b14/B0_39 ;
  wire  \inst_dob_mux_b14/B0_4 ;
  wire  \inst_dob_mux_b14/B0_40 ;
  wire  \inst_dob_mux_b14/B0_41 ;
  wire  \inst_dob_mux_b14/B0_42 ;
  wire  \inst_dob_mux_b14/B0_43 ;
  wire  \inst_dob_mux_b14/B0_44 ;
  wire  \inst_dob_mux_b14/B0_45 ;
  wire  \inst_dob_mux_b14/B0_46 ;
  wire  \inst_dob_mux_b14/B0_47 ;
  wire  \inst_dob_mux_b14/B0_48 ;
  wire  \inst_dob_mux_b14/B0_49 ;
  wire  \inst_dob_mux_b14/B0_5 ;
  wire  \inst_dob_mux_b14/B0_50 ;
  wire  \inst_dob_mux_b14/B0_51 ;
  wire  \inst_dob_mux_b14/B0_52 ;
  wire  \inst_dob_mux_b14/B0_53 ;
  wire  \inst_dob_mux_b14/B0_54 ;
  wire  \inst_dob_mux_b14/B0_55 ;
  wire  \inst_dob_mux_b14/B0_56 ;
  wire  \inst_dob_mux_b14/B0_57 ;
  wire  \inst_dob_mux_b14/B0_58 ;
  wire  \inst_dob_mux_b14/B0_59 ;
  wire  \inst_dob_mux_b14/B0_6 ;
  wire  \inst_dob_mux_b14/B0_60 ;
  wire  \inst_dob_mux_b14/B0_61 ;
  wire  \inst_dob_mux_b14/B0_62 ;
  wire  \inst_dob_mux_b14/B0_63 ;
  wire  \inst_dob_mux_b14/B0_7 ;
  wire  \inst_dob_mux_b14/B0_8 ;
  wire  \inst_dob_mux_b14/B0_9 ;
  wire  \inst_dob_mux_b14/B1_0 ;
  wire  \inst_dob_mux_b14/B1_1 ;
  wire  \inst_dob_mux_b14/B1_10 ;
  wire  \inst_dob_mux_b14/B1_11 ;
  wire  \inst_dob_mux_b14/B1_12 ;
  wire  \inst_dob_mux_b14/B1_13 ;
  wire  \inst_dob_mux_b14/B1_14 ;
  wire  \inst_dob_mux_b14/B1_15 ;
  wire  \inst_dob_mux_b14/B1_16 ;
  wire  \inst_dob_mux_b14/B1_17 ;
  wire  \inst_dob_mux_b14/B1_18 ;
  wire  \inst_dob_mux_b14/B1_19 ;
  wire  \inst_dob_mux_b14/B1_2 ;
  wire  \inst_dob_mux_b14/B1_20 ;
  wire  \inst_dob_mux_b14/B1_21 ;
  wire  \inst_dob_mux_b14/B1_22 ;
  wire  \inst_dob_mux_b14/B1_23 ;
  wire  \inst_dob_mux_b14/B1_24 ;
  wire  \inst_dob_mux_b14/B1_25 ;
  wire  \inst_dob_mux_b14/B1_26 ;
  wire  \inst_dob_mux_b14/B1_27 ;
  wire  \inst_dob_mux_b14/B1_28 ;
  wire  \inst_dob_mux_b14/B1_29 ;
  wire  \inst_dob_mux_b14/B1_3 ;
  wire  \inst_dob_mux_b14/B1_30 ;
  wire  \inst_dob_mux_b14/B1_31 ;
  wire  \inst_dob_mux_b14/B1_4 ;
  wire  \inst_dob_mux_b14/B1_5 ;
  wire  \inst_dob_mux_b14/B1_6 ;
  wire  \inst_dob_mux_b14/B1_7 ;
  wire  \inst_dob_mux_b14/B1_8 ;
  wire  \inst_dob_mux_b14/B1_9 ;
  wire  \inst_dob_mux_b14/B2_0 ;
  wire  \inst_dob_mux_b14/B2_1 ;
  wire  \inst_dob_mux_b14/B2_10 ;
  wire  \inst_dob_mux_b14/B2_11 ;
  wire  \inst_dob_mux_b14/B2_12 ;
  wire  \inst_dob_mux_b14/B2_13 ;
  wire  \inst_dob_mux_b14/B2_14 ;
  wire  \inst_dob_mux_b14/B2_15 ;
  wire  \inst_dob_mux_b14/B2_2 ;
  wire  \inst_dob_mux_b14/B2_3 ;
  wire  \inst_dob_mux_b14/B2_4 ;
  wire  \inst_dob_mux_b14/B2_5 ;
  wire  \inst_dob_mux_b14/B2_6 ;
  wire  \inst_dob_mux_b14/B2_7 ;
  wire  \inst_dob_mux_b14/B2_8 ;
  wire  \inst_dob_mux_b14/B2_9 ;
  wire  \inst_dob_mux_b14/B3_0 ;
  wire  \inst_dob_mux_b14/B3_1 ;
  wire  \inst_dob_mux_b14/B3_2 ;
  wire  \inst_dob_mux_b14/B3_3 ;
  wire  \inst_dob_mux_b14/B3_4 ;
  wire  \inst_dob_mux_b14/B3_5 ;
  wire  \inst_dob_mux_b14/B3_6 ;
  wire  \inst_dob_mux_b14/B3_7 ;
  wire  \inst_dob_mux_b14/B4_0 ;
  wire  \inst_dob_mux_b14/B4_1 ;
  wire  \inst_dob_mux_b14/B4_2 ;
  wire  \inst_dob_mux_b14/B4_3 ;
  wire  \inst_dob_mux_b14/B5_0 ;
  wire  \inst_dob_mux_b14/B5_1 ;
  wire  \inst_dob_mux_b15/B0_0 ;
  wire  \inst_dob_mux_b15/B0_1 ;
  wire  \inst_dob_mux_b15/B0_10 ;
  wire  \inst_dob_mux_b15/B0_11 ;
  wire  \inst_dob_mux_b15/B0_12 ;
  wire  \inst_dob_mux_b15/B0_13 ;
  wire  \inst_dob_mux_b15/B0_14 ;
  wire  \inst_dob_mux_b15/B0_15 ;
  wire  \inst_dob_mux_b15/B0_16 ;
  wire  \inst_dob_mux_b15/B0_17 ;
  wire  \inst_dob_mux_b15/B0_18 ;
  wire  \inst_dob_mux_b15/B0_19 ;
  wire  \inst_dob_mux_b15/B0_2 ;
  wire  \inst_dob_mux_b15/B0_20 ;
  wire  \inst_dob_mux_b15/B0_21 ;
  wire  \inst_dob_mux_b15/B0_22 ;
  wire  \inst_dob_mux_b15/B0_23 ;
  wire  \inst_dob_mux_b15/B0_24 ;
  wire  \inst_dob_mux_b15/B0_25 ;
  wire  \inst_dob_mux_b15/B0_26 ;
  wire  \inst_dob_mux_b15/B0_27 ;
  wire  \inst_dob_mux_b15/B0_28 ;
  wire  \inst_dob_mux_b15/B0_29 ;
  wire  \inst_dob_mux_b15/B0_3 ;
  wire  \inst_dob_mux_b15/B0_30 ;
  wire  \inst_dob_mux_b15/B0_31 ;
  wire  \inst_dob_mux_b15/B0_32 ;
  wire  \inst_dob_mux_b15/B0_33 ;
  wire  \inst_dob_mux_b15/B0_34 ;
  wire  \inst_dob_mux_b15/B0_35 ;
  wire  \inst_dob_mux_b15/B0_36 ;
  wire  \inst_dob_mux_b15/B0_37 ;
  wire  \inst_dob_mux_b15/B0_38 ;
  wire  \inst_dob_mux_b15/B0_39 ;
  wire  \inst_dob_mux_b15/B0_4 ;
  wire  \inst_dob_mux_b15/B0_40 ;
  wire  \inst_dob_mux_b15/B0_41 ;
  wire  \inst_dob_mux_b15/B0_42 ;
  wire  \inst_dob_mux_b15/B0_43 ;
  wire  \inst_dob_mux_b15/B0_44 ;
  wire  \inst_dob_mux_b15/B0_45 ;
  wire  \inst_dob_mux_b15/B0_46 ;
  wire  \inst_dob_mux_b15/B0_47 ;
  wire  \inst_dob_mux_b15/B0_48 ;
  wire  \inst_dob_mux_b15/B0_49 ;
  wire  \inst_dob_mux_b15/B0_5 ;
  wire  \inst_dob_mux_b15/B0_50 ;
  wire  \inst_dob_mux_b15/B0_51 ;
  wire  \inst_dob_mux_b15/B0_52 ;
  wire  \inst_dob_mux_b15/B0_53 ;
  wire  \inst_dob_mux_b15/B0_54 ;
  wire  \inst_dob_mux_b15/B0_55 ;
  wire  \inst_dob_mux_b15/B0_56 ;
  wire  \inst_dob_mux_b15/B0_57 ;
  wire  \inst_dob_mux_b15/B0_58 ;
  wire  \inst_dob_mux_b15/B0_59 ;
  wire  \inst_dob_mux_b15/B0_6 ;
  wire  \inst_dob_mux_b15/B0_60 ;
  wire  \inst_dob_mux_b15/B0_61 ;
  wire  \inst_dob_mux_b15/B0_62 ;
  wire  \inst_dob_mux_b15/B0_63 ;
  wire  \inst_dob_mux_b15/B0_7 ;
  wire  \inst_dob_mux_b15/B0_8 ;
  wire  \inst_dob_mux_b15/B0_9 ;
  wire  \inst_dob_mux_b15/B1_0 ;
  wire  \inst_dob_mux_b15/B1_1 ;
  wire  \inst_dob_mux_b15/B1_10 ;
  wire  \inst_dob_mux_b15/B1_11 ;
  wire  \inst_dob_mux_b15/B1_12 ;
  wire  \inst_dob_mux_b15/B1_13 ;
  wire  \inst_dob_mux_b15/B1_14 ;
  wire  \inst_dob_mux_b15/B1_15 ;
  wire  \inst_dob_mux_b15/B1_16 ;
  wire  \inst_dob_mux_b15/B1_17 ;
  wire  \inst_dob_mux_b15/B1_18 ;
  wire  \inst_dob_mux_b15/B1_19 ;
  wire  \inst_dob_mux_b15/B1_2 ;
  wire  \inst_dob_mux_b15/B1_20 ;
  wire  \inst_dob_mux_b15/B1_21 ;
  wire  \inst_dob_mux_b15/B1_22 ;
  wire  \inst_dob_mux_b15/B1_23 ;
  wire  \inst_dob_mux_b15/B1_24 ;
  wire  \inst_dob_mux_b15/B1_25 ;
  wire  \inst_dob_mux_b15/B1_26 ;
  wire  \inst_dob_mux_b15/B1_27 ;
  wire  \inst_dob_mux_b15/B1_28 ;
  wire  \inst_dob_mux_b15/B1_29 ;
  wire  \inst_dob_mux_b15/B1_3 ;
  wire  \inst_dob_mux_b15/B1_30 ;
  wire  \inst_dob_mux_b15/B1_31 ;
  wire  \inst_dob_mux_b15/B1_4 ;
  wire  \inst_dob_mux_b15/B1_5 ;
  wire  \inst_dob_mux_b15/B1_6 ;
  wire  \inst_dob_mux_b15/B1_7 ;
  wire  \inst_dob_mux_b15/B1_8 ;
  wire  \inst_dob_mux_b15/B1_9 ;
  wire  \inst_dob_mux_b15/B2_0 ;
  wire  \inst_dob_mux_b15/B2_1 ;
  wire  \inst_dob_mux_b15/B2_10 ;
  wire  \inst_dob_mux_b15/B2_11 ;
  wire  \inst_dob_mux_b15/B2_12 ;
  wire  \inst_dob_mux_b15/B2_13 ;
  wire  \inst_dob_mux_b15/B2_14 ;
  wire  \inst_dob_mux_b15/B2_15 ;
  wire  \inst_dob_mux_b15/B2_2 ;
  wire  \inst_dob_mux_b15/B2_3 ;
  wire  \inst_dob_mux_b15/B2_4 ;
  wire  \inst_dob_mux_b15/B2_5 ;
  wire  \inst_dob_mux_b15/B2_6 ;
  wire  \inst_dob_mux_b15/B2_7 ;
  wire  \inst_dob_mux_b15/B2_8 ;
  wire  \inst_dob_mux_b15/B2_9 ;
  wire  \inst_dob_mux_b15/B3_0 ;
  wire  \inst_dob_mux_b15/B3_1 ;
  wire  \inst_dob_mux_b15/B3_2 ;
  wire  \inst_dob_mux_b15/B3_3 ;
  wire  \inst_dob_mux_b15/B3_4 ;
  wire  \inst_dob_mux_b15/B3_5 ;
  wire  \inst_dob_mux_b15/B3_6 ;
  wire  \inst_dob_mux_b15/B3_7 ;
  wire  \inst_dob_mux_b15/B4_0 ;
  wire  \inst_dob_mux_b15/B4_1 ;
  wire  \inst_dob_mux_b15/B4_2 ;
  wire  \inst_dob_mux_b15/B4_3 ;
  wire  \inst_dob_mux_b15/B5_0 ;
  wire  \inst_dob_mux_b15/B5_1 ;
  wire  \inst_dob_mux_b2/B0_0 ;
  wire  \inst_dob_mux_b2/B0_1 ;
  wire  \inst_dob_mux_b2/B0_10 ;
  wire  \inst_dob_mux_b2/B0_11 ;
  wire  \inst_dob_mux_b2/B0_12 ;
  wire  \inst_dob_mux_b2/B0_13 ;
  wire  \inst_dob_mux_b2/B0_14 ;
  wire  \inst_dob_mux_b2/B0_15 ;
  wire  \inst_dob_mux_b2/B0_16 ;
  wire  \inst_dob_mux_b2/B0_17 ;
  wire  \inst_dob_mux_b2/B0_18 ;
  wire  \inst_dob_mux_b2/B0_19 ;
  wire  \inst_dob_mux_b2/B0_2 ;
  wire  \inst_dob_mux_b2/B0_20 ;
  wire  \inst_dob_mux_b2/B0_21 ;
  wire  \inst_dob_mux_b2/B0_22 ;
  wire  \inst_dob_mux_b2/B0_23 ;
  wire  \inst_dob_mux_b2/B0_24 ;
  wire  \inst_dob_mux_b2/B0_25 ;
  wire  \inst_dob_mux_b2/B0_26 ;
  wire  \inst_dob_mux_b2/B0_27 ;
  wire  \inst_dob_mux_b2/B0_28 ;
  wire  \inst_dob_mux_b2/B0_29 ;
  wire  \inst_dob_mux_b2/B0_3 ;
  wire  \inst_dob_mux_b2/B0_30 ;
  wire  \inst_dob_mux_b2/B0_31 ;
  wire  \inst_dob_mux_b2/B0_32 ;
  wire  \inst_dob_mux_b2/B0_33 ;
  wire  \inst_dob_mux_b2/B0_34 ;
  wire  \inst_dob_mux_b2/B0_35 ;
  wire  \inst_dob_mux_b2/B0_36 ;
  wire  \inst_dob_mux_b2/B0_37 ;
  wire  \inst_dob_mux_b2/B0_38 ;
  wire  \inst_dob_mux_b2/B0_39 ;
  wire  \inst_dob_mux_b2/B0_4 ;
  wire  \inst_dob_mux_b2/B0_40 ;
  wire  \inst_dob_mux_b2/B0_41 ;
  wire  \inst_dob_mux_b2/B0_42 ;
  wire  \inst_dob_mux_b2/B0_43 ;
  wire  \inst_dob_mux_b2/B0_44 ;
  wire  \inst_dob_mux_b2/B0_45 ;
  wire  \inst_dob_mux_b2/B0_46 ;
  wire  \inst_dob_mux_b2/B0_47 ;
  wire  \inst_dob_mux_b2/B0_48 ;
  wire  \inst_dob_mux_b2/B0_49 ;
  wire  \inst_dob_mux_b2/B0_5 ;
  wire  \inst_dob_mux_b2/B0_50 ;
  wire  \inst_dob_mux_b2/B0_51 ;
  wire  \inst_dob_mux_b2/B0_52 ;
  wire  \inst_dob_mux_b2/B0_53 ;
  wire  \inst_dob_mux_b2/B0_54 ;
  wire  \inst_dob_mux_b2/B0_55 ;
  wire  \inst_dob_mux_b2/B0_56 ;
  wire  \inst_dob_mux_b2/B0_57 ;
  wire  \inst_dob_mux_b2/B0_58 ;
  wire  \inst_dob_mux_b2/B0_59 ;
  wire  \inst_dob_mux_b2/B0_6 ;
  wire  \inst_dob_mux_b2/B0_60 ;
  wire  \inst_dob_mux_b2/B0_61 ;
  wire  \inst_dob_mux_b2/B0_62 ;
  wire  \inst_dob_mux_b2/B0_63 ;
  wire  \inst_dob_mux_b2/B0_7 ;
  wire  \inst_dob_mux_b2/B0_8 ;
  wire  \inst_dob_mux_b2/B0_9 ;
  wire  \inst_dob_mux_b2/B1_0 ;
  wire  \inst_dob_mux_b2/B1_1 ;
  wire  \inst_dob_mux_b2/B1_10 ;
  wire  \inst_dob_mux_b2/B1_11 ;
  wire  \inst_dob_mux_b2/B1_12 ;
  wire  \inst_dob_mux_b2/B1_13 ;
  wire  \inst_dob_mux_b2/B1_14 ;
  wire  \inst_dob_mux_b2/B1_15 ;
  wire  \inst_dob_mux_b2/B1_16 ;
  wire  \inst_dob_mux_b2/B1_17 ;
  wire  \inst_dob_mux_b2/B1_18 ;
  wire  \inst_dob_mux_b2/B1_19 ;
  wire  \inst_dob_mux_b2/B1_2 ;
  wire  \inst_dob_mux_b2/B1_20 ;
  wire  \inst_dob_mux_b2/B1_21 ;
  wire  \inst_dob_mux_b2/B1_22 ;
  wire  \inst_dob_mux_b2/B1_23 ;
  wire  \inst_dob_mux_b2/B1_24 ;
  wire  \inst_dob_mux_b2/B1_25 ;
  wire  \inst_dob_mux_b2/B1_26 ;
  wire  \inst_dob_mux_b2/B1_27 ;
  wire  \inst_dob_mux_b2/B1_28 ;
  wire  \inst_dob_mux_b2/B1_29 ;
  wire  \inst_dob_mux_b2/B1_3 ;
  wire  \inst_dob_mux_b2/B1_30 ;
  wire  \inst_dob_mux_b2/B1_31 ;
  wire  \inst_dob_mux_b2/B1_4 ;
  wire  \inst_dob_mux_b2/B1_5 ;
  wire  \inst_dob_mux_b2/B1_6 ;
  wire  \inst_dob_mux_b2/B1_7 ;
  wire  \inst_dob_mux_b2/B1_8 ;
  wire  \inst_dob_mux_b2/B1_9 ;
  wire  \inst_dob_mux_b2/B2_0 ;
  wire  \inst_dob_mux_b2/B2_1 ;
  wire  \inst_dob_mux_b2/B2_10 ;
  wire  \inst_dob_mux_b2/B2_11 ;
  wire  \inst_dob_mux_b2/B2_12 ;
  wire  \inst_dob_mux_b2/B2_13 ;
  wire  \inst_dob_mux_b2/B2_14 ;
  wire  \inst_dob_mux_b2/B2_15 ;
  wire  \inst_dob_mux_b2/B2_2 ;
  wire  \inst_dob_mux_b2/B2_3 ;
  wire  \inst_dob_mux_b2/B2_4 ;
  wire  \inst_dob_mux_b2/B2_5 ;
  wire  \inst_dob_mux_b2/B2_6 ;
  wire  \inst_dob_mux_b2/B2_7 ;
  wire  \inst_dob_mux_b2/B2_8 ;
  wire  \inst_dob_mux_b2/B2_9 ;
  wire  \inst_dob_mux_b2/B3_0 ;
  wire  \inst_dob_mux_b2/B3_1 ;
  wire  \inst_dob_mux_b2/B3_2 ;
  wire  \inst_dob_mux_b2/B3_3 ;
  wire  \inst_dob_mux_b2/B3_4 ;
  wire  \inst_dob_mux_b2/B3_5 ;
  wire  \inst_dob_mux_b2/B3_6 ;
  wire  \inst_dob_mux_b2/B3_7 ;
  wire  \inst_dob_mux_b2/B4_0 ;
  wire  \inst_dob_mux_b2/B4_1 ;
  wire  \inst_dob_mux_b2/B4_2 ;
  wire  \inst_dob_mux_b2/B4_3 ;
  wire  \inst_dob_mux_b2/B5_0 ;
  wire  \inst_dob_mux_b2/B5_1 ;
  wire  \inst_dob_mux_b3/B0_0 ;
  wire  \inst_dob_mux_b3/B0_1 ;
  wire  \inst_dob_mux_b3/B0_10 ;
  wire  \inst_dob_mux_b3/B0_11 ;
  wire  \inst_dob_mux_b3/B0_12 ;
  wire  \inst_dob_mux_b3/B0_13 ;
  wire  \inst_dob_mux_b3/B0_14 ;
  wire  \inst_dob_mux_b3/B0_15 ;
  wire  \inst_dob_mux_b3/B0_16 ;
  wire  \inst_dob_mux_b3/B0_17 ;
  wire  \inst_dob_mux_b3/B0_18 ;
  wire  \inst_dob_mux_b3/B0_19 ;
  wire  \inst_dob_mux_b3/B0_2 ;
  wire  \inst_dob_mux_b3/B0_20 ;
  wire  \inst_dob_mux_b3/B0_21 ;
  wire  \inst_dob_mux_b3/B0_22 ;
  wire  \inst_dob_mux_b3/B0_23 ;
  wire  \inst_dob_mux_b3/B0_24 ;
  wire  \inst_dob_mux_b3/B0_25 ;
  wire  \inst_dob_mux_b3/B0_26 ;
  wire  \inst_dob_mux_b3/B0_27 ;
  wire  \inst_dob_mux_b3/B0_28 ;
  wire  \inst_dob_mux_b3/B0_29 ;
  wire  \inst_dob_mux_b3/B0_3 ;
  wire  \inst_dob_mux_b3/B0_30 ;
  wire  \inst_dob_mux_b3/B0_31 ;
  wire  \inst_dob_mux_b3/B0_32 ;
  wire  \inst_dob_mux_b3/B0_33 ;
  wire  \inst_dob_mux_b3/B0_34 ;
  wire  \inst_dob_mux_b3/B0_35 ;
  wire  \inst_dob_mux_b3/B0_36 ;
  wire  \inst_dob_mux_b3/B0_37 ;
  wire  \inst_dob_mux_b3/B0_38 ;
  wire  \inst_dob_mux_b3/B0_39 ;
  wire  \inst_dob_mux_b3/B0_4 ;
  wire  \inst_dob_mux_b3/B0_40 ;
  wire  \inst_dob_mux_b3/B0_41 ;
  wire  \inst_dob_mux_b3/B0_42 ;
  wire  \inst_dob_mux_b3/B0_43 ;
  wire  \inst_dob_mux_b3/B0_44 ;
  wire  \inst_dob_mux_b3/B0_45 ;
  wire  \inst_dob_mux_b3/B0_46 ;
  wire  \inst_dob_mux_b3/B0_47 ;
  wire  \inst_dob_mux_b3/B0_48 ;
  wire  \inst_dob_mux_b3/B0_49 ;
  wire  \inst_dob_mux_b3/B0_5 ;
  wire  \inst_dob_mux_b3/B0_50 ;
  wire  \inst_dob_mux_b3/B0_51 ;
  wire  \inst_dob_mux_b3/B0_52 ;
  wire  \inst_dob_mux_b3/B0_53 ;
  wire  \inst_dob_mux_b3/B0_54 ;
  wire  \inst_dob_mux_b3/B0_55 ;
  wire  \inst_dob_mux_b3/B0_56 ;
  wire  \inst_dob_mux_b3/B0_57 ;
  wire  \inst_dob_mux_b3/B0_58 ;
  wire  \inst_dob_mux_b3/B0_59 ;
  wire  \inst_dob_mux_b3/B0_6 ;
  wire  \inst_dob_mux_b3/B0_60 ;
  wire  \inst_dob_mux_b3/B0_61 ;
  wire  \inst_dob_mux_b3/B0_62 ;
  wire  \inst_dob_mux_b3/B0_63 ;
  wire  \inst_dob_mux_b3/B0_7 ;
  wire  \inst_dob_mux_b3/B0_8 ;
  wire  \inst_dob_mux_b3/B0_9 ;
  wire  \inst_dob_mux_b3/B1_0 ;
  wire  \inst_dob_mux_b3/B1_1 ;
  wire  \inst_dob_mux_b3/B1_10 ;
  wire  \inst_dob_mux_b3/B1_11 ;
  wire  \inst_dob_mux_b3/B1_12 ;
  wire  \inst_dob_mux_b3/B1_13 ;
  wire  \inst_dob_mux_b3/B1_14 ;
  wire  \inst_dob_mux_b3/B1_15 ;
  wire  \inst_dob_mux_b3/B1_16 ;
  wire  \inst_dob_mux_b3/B1_17 ;
  wire  \inst_dob_mux_b3/B1_18 ;
  wire  \inst_dob_mux_b3/B1_19 ;
  wire  \inst_dob_mux_b3/B1_2 ;
  wire  \inst_dob_mux_b3/B1_20 ;
  wire  \inst_dob_mux_b3/B1_21 ;
  wire  \inst_dob_mux_b3/B1_22 ;
  wire  \inst_dob_mux_b3/B1_23 ;
  wire  \inst_dob_mux_b3/B1_24 ;
  wire  \inst_dob_mux_b3/B1_25 ;
  wire  \inst_dob_mux_b3/B1_26 ;
  wire  \inst_dob_mux_b3/B1_27 ;
  wire  \inst_dob_mux_b3/B1_28 ;
  wire  \inst_dob_mux_b3/B1_29 ;
  wire  \inst_dob_mux_b3/B1_3 ;
  wire  \inst_dob_mux_b3/B1_30 ;
  wire  \inst_dob_mux_b3/B1_31 ;
  wire  \inst_dob_mux_b3/B1_4 ;
  wire  \inst_dob_mux_b3/B1_5 ;
  wire  \inst_dob_mux_b3/B1_6 ;
  wire  \inst_dob_mux_b3/B1_7 ;
  wire  \inst_dob_mux_b3/B1_8 ;
  wire  \inst_dob_mux_b3/B1_9 ;
  wire  \inst_dob_mux_b3/B2_0 ;
  wire  \inst_dob_mux_b3/B2_1 ;
  wire  \inst_dob_mux_b3/B2_10 ;
  wire  \inst_dob_mux_b3/B2_11 ;
  wire  \inst_dob_mux_b3/B2_12 ;
  wire  \inst_dob_mux_b3/B2_13 ;
  wire  \inst_dob_mux_b3/B2_14 ;
  wire  \inst_dob_mux_b3/B2_15 ;
  wire  \inst_dob_mux_b3/B2_2 ;
  wire  \inst_dob_mux_b3/B2_3 ;
  wire  \inst_dob_mux_b3/B2_4 ;
  wire  \inst_dob_mux_b3/B2_5 ;
  wire  \inst_dob_mux_b3/B2_6 ;
  wire  \inst_dob_mux_b3/B2_7 ;
  wire  \inst_dob_mux_b3/B2_8 ;
  wire  \inst_dob_mux_b3/B2_9 ;
  wire  \inst_dob_mux_b3/B3_0 ;
  wire  \inst_dob_mux_b3/B3_1 ;
  wire  \inst_dob_mux_b3/B3_2 ;
  wire  \inst_dob_mux_b3/B3_3 ;
  wire  \inst_dob_mux_b3/B3_4 ;
  wire  \inst_dob_mux_b3/B3_5 ;
  wire  \inst_dob_mux_b3/B3_6 ;
  wire  \inst_dob_mux_b3/B3_7 ;
  wire  \inst_dob_mux_b3/B4_0 ;
  wire  \inst_dob_mux_b3/B4_1 ;
  wire  \inst_dob_mux_b3/B4_2 ;
  wire  \inst_dob_mux_b3/B4_3 ;
  wire  \inst_dob_mux_b3/B5_0 ;
  wire  \inst_dob_mux_b3/B5_1 ;
  wire  \inst_dob_mux_b4/B0_0 ;
  wire  \inst_dob_mux_b4/B0_1 ;
  wire  \inst_dob_mux_b4/B0_10 ;
  wire  \inst_dob_mux_b4/B0_11 ;
  wire  \inst_dob_mux_b4/B0_12 ;
  wire  \inst_dob_mux_b4/B0_13 ;
  wire  \inst_dob_mux_b4/B0_14 ;
  wire  \inst_dob_mux_b4/B0_15 ;
  wire  \inst_dob_mux_b4/B0_16 ;
  wire  \inst_dob_mux_b4/B0_17 ;
  wire  \inst_dob_mux_b4/B0_18 ;
  wire  \inst_dob_mux_b4/B0_19 ;
  wire  \inst_dob_mux_b4/B0_2 ;
  wire  \inst_dob_mux_b4/B0_20 ;
  wire  \inst_dob_mux_b4/B0_21 ;
  wire  \inst_dob_mux_b4/B0_22 ;
  wire  \inst_dob_mux_b4/B0_23 ;
  wire  \inst_dob_mux_b4/B0_24 ;
  wire  \inst_dob_mux_b4/B0_25 ;
  wire  \inst_dob_mux_b4/B0_26 ;
  wire  \inst_dob_mux_b4/B0_27 ;
  wire  \inst_dob_mux_b4/B0_28 ;
  wire  \inst_dob_mux_b4/B0_29 ;
  wire  \inst_dob_mux_b4/B0_3 ;
  wire  \inst_dob_mux_b4/B0_30 ;
  wire  \inst_dob_mux_b4/B0_31 ;
  wire  \inst_dob_mux_b4/B0_32 ;
  wire  \inst_dob_mux_b4/B0_33 ;
  wire  \inst_dob_mux_b4/B0_34 ;
  wire  \inst_dob_mux_b4/B0_35 ;
  wire  \inst_dob_mux_b4/B0_36 ;
  wire  \inst_dob_mux_b4/B0_37 ;
  wire  \inst_dob_mux_b4/B0_38 ;
  wire  \inst_dob_mux_b4/B0_39 ;
  wire  \inst_dob_mux_b4/B0_4 ;
  wire  \inst_dob_mux_b4/B0_40 ;
  wire  \inst_dob_mux_b4/B0_41 ;
  wire  \inst_dob_mux_b4/B0_42 ;
  wire  \inst_dob_mux_b4/B0_43 ;
  wire  \inst_dob_mux_b4/B0_44 ;
  wire  \inst_dob_mux_b4/B0_45 ;
  wire  \inst_dob_mux_b4/B0_46 ;
  wire  \inst_dob_mux_b4/B0_47 ;
  wire  \inst_dob_mux_b4/B0_48 ;
  wire  \inst_dob_mux_b4/B0_49 ;
  wire  \inst_dob_mux_b4/B0_5 ;
  wire  \inst_dob_mux_b4/B0_50 ;
  wire  \inst_dob_mux_b4/B0_51 ;
  wire  \inst_dob_mux_b4/B0_52 ;
  wire  \inst_dob_mux_b4/B0_53 ;
  wire  \inst_dob_mux_b4/B0_54 ;
  wire  \inst_dob_mux_b4/B0_55 ;
  wire  \inst_dob_mux_b4/B0_56 ;
  wire  \inst_dob_mux_b4/B0_57 ;
  wire  \inst_dob_mux_b4/B0_58 ;
  wire  \inst_dob_mux_b4/B0_59 ;
  wire  \inst_dob_mux_b4/B0_6 ;
  wire  \inst_dob_mux_b4/B0_60 ;
  wire  \inst_dob_mux_b4/B0_61 ;
  wire  \inst_dob_mux_b4/B0_62 ;
  wire  \inst_dob_mux_b4/B0_63 ;
  wire  \inst_dob_mux_b4/B0_7 ;
  wire  \inst_dob_mux_b4/B0_8 ;
  wire  \inst_dob_mux_b4/B0_9 ;
  wire  \inst_dob_mux_b4/B1_0 ;
  wire  \inst_dob_mux_b4/B1_1 ;
  wire  \inst_dob_mux_b4/B1_10 ;
  wire  \inst_dob_mux_b4/B1_11 ;
  wire  \inst_dob_mux_b4/B1_12 ;
  wire  \inst_dob_mux_b4/B1_13 ;
  wire  \inst_dob_mux_b4/B1_14 ;
  wire  \inst_dob_mux_b4/B1_15 ;
  wire  \inst_dob_mux_b4/B1_16 ;
  wire  \inst_dob_mux_b4/B1_17 ;
  wire  \inst_dob_mux_b4/B1_18 ;
  wire  \inst_dob_mux_b4/B1_19 ;
  wire  \inst_dob_mux_b4/B1_2 ;
  wire  \inst_dob_mux_b4/B1_20 ;
  wire  \inst_dob_mux_b4/B1_21 ;
  wire  \inst_dob_mux_b4/B1_22 ;
  wire  \inst_dob_mux_b4/B1_23 ;
  wire  \inst_dob_mux_b4/B1_24 ;
  wire  \inst_dob_mux_b4/B1_25 ;
  wire  \inst_dob_mux_b4/B1_26 ;
  wire  \inst_dob_mux_b4/B1_27 ;
  wire  \inst_dob_mux_b4/B1_28 ;
  wire  \inst_dob_mux_b4/B1_29 ;
  wire  \inst_dob_mux_b4/B1_3 ;
  wire  \inst_dob_mux_b4/B1_30 ;
  wire  \inst_dob_mux_b4/B1_31 ;
  wire  \inst_dob_mux_b4/B1_4 ;
  wire  \inst_dob_mux_b4/B1_5 ;
  wire  \inst_dob_mux_b4/B1_6 ;
  wire  \inst_dob_mux_b4/B1_7 ;
  wire  \inst_dob_mux_b4/B1_8 ;
  wire  \inst_dob_mux_b4/B1_9 ;
  wire  \inst_dob_mux_b4/B2_0 ;
  wire  \inst_dob_mux_b4/B2_1 ;
  wire  \inst_dob_mux_b4/B2_10 ;
  wire  \inst_dob_mux_b4/B2_11 ;
  wire  \inst_dob_mux_b4/B2_12 ;
  wire  \inst_dob_mux_b4/B2_13 ;
  wire  \inst_dob_mux_b4/B2_14 ;
  wire  \inst_dob_mux_b4/B2_15 ;
  wire  \inst_dob_mux_b4/B2_2 ;
  wire  \inst_dob_mux_b4/B2_3 ;
  wire  \inst_dob_mux_b4/B2_4 ;
  wire  \inst_dob_mux_b4/B2_5 ;
  wire  \inst_dob_mux_b4/B2_6 ;
  wire  \inst_dob_mux_b4/B2_7 ;
  wire  \inst_dob_mux_b4/B2_8 ;
  wire  \inst_dob_mux_b4/B2_9 ;
  wire  \inst_dob_mux_b4/B3_0 ;
  wire  \inst_dob_mux_b4/B3_1 ;
  wire  \inst_dob_mux_b4/B3_2 ;
  wire  \inst_dob_mux_b4/B3_3 ;
  wire  \inst_dob_mux_b4/B3_4 ;
  wire  \inst_dob_mux_b4/B3_5 ;
  wire  \inst_dob_mux_b4/B3_6 ;
  wire  \inst_dob_mux_b4/B3_7 ;
  wire  \inst_dob_mux_b4/B4_0 ;
  wire  \inst_dob_mux_b4/B4_1 ;
  wire  \inst_dob_mux_b4/B4_2 ;
  wire  \inst_dob_mux_b4/B4_3 ;
  wire  \inst_dob_mux_b4/B5_0 ;
  wire  \inst_dob_mux_b4/B5_1 ;
  wire  \inst_dob_mux_b5/B0_0 ;
  wire  \inst_dob_mux_b5/B0_1 ;
  wire  \inst_dob_mux_b5/B0_10 ;
  wire  \inst_dob_mux_b5/B0_11 ;
  wire  \inst_dob_mux_b5/B0_12 ;
  wire  \inst_dob_mux_b5/B0_13 ;
  wire  \inst_dob_mux_b5/B0_14 ;
  wire  \inst_dob_mux_b5/B0_15 ;
  wire  \inst_dob_mux_b5/B0_16 ;
  wire  \inst_dob_mux_b5/B0_17 ;
  wire  \inst_dob_mux_b5/B0_18 ;
  wire  \inst_dob_mux_b5/B0_19 ;
  wire  \inst_dob_mux_b5/B0_2 ;
  wire  \inst_dob_mux_b5/B0_20 ;
  wire  \inst_dob_mux_b5/B0_21 ;
  wire  \inst_dob_mux_b5/B0_22 ;
  wire  \inst_dob_mux_b5/B0_23 ;
  wire  \inst_dob_mux_b5/B0_24 ;
  wire  \inst_dob_mux_b5/B0_25 ;
  wire  \inst_dob_mux_b5/B0_26 ;
  wire  \inst_dob_mux_b5/B0_27 ;
  wire  \inst_dob_mux_b5/B0_28 ;
  wire  \inst_dob_mux_b5/B0_29 ;
  wire  \inst_dob_mux_b5/B0_3 ;
  wire  \inst_dob_mux_b5/B0_30 ;
  wire  \inst_dob_mux_b5/B0_31 ;
  wire  \inst_dob_mux_b5/B0_32 ;
  wire  \inst_dob_mux_b5/B0_33 ;
  wire  \inst_dob_mux_b5/B0_34 ;
  wire  \inst_dob_mux_b5/B0_35 ;
  wire  \inst_dob_mux_b5/B0_36 ;
  wire  \inst_dob_mux_b5/B0_37 ;
  wire  \inst_dob_mux_b5/B0_38 ;
  wire  \inst_dob_mux_b5/B0_39 ;
  wire  \inst_dob_mux_b5/B0_4 ;
  wire  \inst_dob_mux_b5/B0_40 ;
  wire  \inst_dob_mux_b5/B0_41 ;
  wire  \inst_dob_mux_b5/B0_42 ;
  wire  \inst_dob_mux_b5/B0_43 ;
  wire  \inst_dob_mux_b5/B0_44 ;
  wire  \inst_dob_mux_b5/B0_45 ;
  wire  \inst_dob_mux_b5/B0_46 ;
  wire  \inst_dob_mux_b5/B0_47 ;
  wire  \inst_dob_mux_b5/B0_48 ;
  wire  \inst_dob_mux_b5/B0_49 ;
  wire  \inst_dob_mux_b5/B0_5 ;
  wire  \inst_dob_mux_b5/B0_50 ;
  wire  \inst_dob_mux_b5/B0_51 ;
  wire  \inst_dob_mux_b5/B0_52 ;
  wire  \inst_dob_mux_b5/B0_53 ;
  wire  \inst_dob_mux_b5/B0_54 ;
  wire  \inst_dob_mux_b5/B0_55 ;
  wire  \inst_dob_mux_b5/B0_56 ;
  wire  \inst_dob_mux_b5/B0_57 ;
  wire  \inst_dob_mux_b5/B0_58 ;
  wire  \inst_dob_mux_b5/B0_59 ;
  wire  \inst_dob_mux_b5/B0_6 ;
  wire  \inst_dob_mux_b5/B0_60 ;
  wire  \inst_dob_mux_b5/B0_61 ;
  wire  \inst_dob_mux_b5/B0_62 ;
  wire  \inst_dob_mux_b5/B0_63 ;
  wire  \inst_dob_mux_b5/B0_7 ;
  wire  \inst_dob_mux_b5/B0_8 ;
  wire  \inst_dob_mux_b5/B0_9 ;
  wire  \inst_dob_mux_b5/B1_0 ;
  wire  \inst_dob_mux_b5/B1_1 ;
  wire  \inst_dob_mux_b5/B1_10 ;
  wire  \inst_dob_mux_b5/B1_11 ;
  wire  \inst_dob_mux_b5/B1_12 ;
  wire  \inst_dob_mux_b5/B1_13 ;
  wire  \inst_dob_mux_b5/B1_14 ;
  wire  \inst_dob_mux_b5/B1_15 ;
  wire  \inst_dob_mux_b5/B1_16 ;
  wire  \inst_dob_mux_b5/B1_17 ;
  wire  \inst_dob_mux_b5/B1_18 ;
  wire  \inst_dob_mux_b5/B1_19 ;
  wire  \inst_dob_mux_b5/B1_2 ;
  wire  \inst_dob_mux_b5/B1_20 ;
  wire  \inst_dob_mux_b5/B1_21 ;
  wire  \inst_dob_mux_b5/B1_22 ;
  wire  \inst_dob_mux_b5/B1_23 ;
  wire  \inst_dob_mux_b5/B1_24 ;
  wire  \inst_dob_mux_b5/B1_25 ;
  wire  \inst_dob_mux_b5/B1_26 ;
  wire  \inst_dob_mux_b5/B1_27 ;
  wire  \inst_dob_mux_b5/B1_28 ;
  wire  \inst_dob_mux_b5/B1_29 ;
  wire  \inst_dob_mux_b5/B1_3 ;
  wire  \inst_dob_mux_b5/B1_30 ;
  wire  \inst_dob_mux_b5/B1_31 ;
  wire  \inst_dob_mux_b5/B1_4 ;
  wire  \inst_dob_mux_b5/B1_5 ;
  wire  \inst_dob_mux_b5/B1_6 ;
  wire  \inst_dob_mux_b5/B1_7 ;
  wire  \inst_dob_mux_b5/B1_8 ;
  wire  \inst_dob_mux_b5/B1_9 ;
  wire  \inst_dob_mux_b5/B2_0 ;
  wire  \inst_dob_mux_b5/B2_1 ;
  wire  \inst_dob_mux_b5/B2_10 ;
  wire  \inst_dob_mux_b5/B2_11 ;
  wire  \inst_dob_mux_b5/B2_12 ;
  wire  \inst_dob_mux_b5/B2_13 ;
  wire  \inst_dob_mux_b5/B2_14 ;
  wire  \inst_dob_mux_b5/B2_15 ;
  wire  \inst_dob_mux_b5/B2_2 ;
  wire  \inst_dob_mux_b5/B2_3 ;
  wire  \inst_dob_mux_b5/B2_4 ;
  wire  \inst_dob_mux_b5/B2_5 ;
  wire  \inst_dob_mux_b5/B2_6 ;
  wire  \inst_dob_mux_b5/B2_7 ;
  wire  \inst_dob_mux_b5/B2_8 ;
  wire  \inst_dob_mux_b5/B2_9 ;
  wire  \inst_dob_mux_b5/B3_0 ;
  wire  \inst_dob_mux_b5/B3_1 ;
  wire  \inst_dob_mux_b5/B3_2 ;
  wire  \inst_dob_mux_b5/B3_3 ;
  wire  \inst_dob_mux_b5/B3_4 ;
  wire  \inst_dob_mux_b5/B3_5 ;
  wire  \inst_dob_mux_b5/B3_6 ;
  wire  \inst_dob_mux_b5/B3_7 ;
  wire  \inst_dob_mux_b5/B4_0 ;
  wire  \inst_dob_mux_b5/B4_1 ;
  wire  \inst_dob_mux_b5/B4_2 ;
  wire  \inst_dob_mux_b5/B4_3 ;
  wire  \inst_dob_mux_b5/B5_0 ;
  wire  \inst_dob_mux_b5/B5_1 ;
  wire  \inst_dob_mux_b6/B0_0 ;
  wire  \inst_dob_mux_b6/B0_1 ;
  wire  \inst_dob_mux_b6/B0_10 ;
  wire  \inst_dob_mux_b6/B0_11 ;
  wire  \inst_dob_mux_b6/B0_12 ;
  wire  \inst_dob_mux_b6/B0_13 ;
  wire  \inst_dob_mux_b6/B0_14 ;
  wire  \inst_dob_mux_b6/B0_15 ;
  wire  \inst_dob_mux_b6/B0_16 ;
  wire  \inst_dob_mux_b6/B0_17 ;
  wire  \inst_dob_mux_b6/B0_18 ;
  wire  \inst_dob_mux_b6/B0_19 ;
  wire  \inst_dob_mux_b6/B0_2 ;
  wire  \inst_dob_mux_b6/B0_20 ;
  wire  \inst_dob_mux_b6/B0_21 ;
  wire  \inst_dob_mux_b6/B0_22 ;
  wire  \inst_dob_mux_b6/B0_23 ;
  wire  \inst_dob_mux_b6/B0_24 ;
  wire  \inst_dob_mux_b6/B0_25 ;
  wire  \inst_dob_mux_b6/B0_26 ;
  wire  \inst_dob_mux_b6/B0_27 ;
  wire  \inst_dob_mux_b6/B0_28 ;
  wire  \inst_dob_mux_b6/B0_29 ;
  wire  \inst_dob_mux_b6/B0_3 ;
  wire  \inst_dob_mux_b6/B0_30 ;
  wire  \inst_dob_mux_b6/B0_31 ;
  wire  \inst_dob_mux_b6/B0_32 ;
  wire  \inst_dob_mux_b6/B0_33 ;
  wire  \inst_dob_mux_b6/B0_34 ;
  wire  \inst_dob_mux_b6/B0_35 ;
  wire  \inst_dob_mux_b6/B0_36 ;
  wire  \inst_dob_mux_b6/B0_37 ;
  wire  \inst_dob_mux_b6/B0_38 ;
  wire  \inst_dob_mux_b6/B0_39 ;
  wire  \inst_dob_mux_b6/B0_4 ;
  wire  \inst_dob_mux_b6/B0_40 ;
  wire  \inst_dob_mux_b6/B0_41 ;
  wire  \inst_dob_mux_b6/B0_42 ;
  wire  \inst_dob_mux_b6/B0_43 ;
  wire  \inst_dob_mux_b6/B0_44 ;
  wire  \inst_dob_mux_b6/B0_45 ;
  wire  \inst_dob_mux_b6/B0_46 ;
  wire  \inst_dob_mux_b6/B0_47 ;
  wire  \inst_dob_mux_b6/B0_48 ;
  wire  \inst_dob_mux_b6/B0_49 ;
  wire  \inst_dob_mux_b6/B0_5 ;
  wire  \inst_dob_mux_b6/B0_50 ;
  wire  \inst_dob_mux_b6/B0_51 ;
  wire  \inst_dob_mux_b6/B0_52 ;
  wire  \inst_dob_mux_b6/B0_53 ;
  wire  \inst_dob_mux_b6/B0_54 ;
  wire  \inst_dob_mux_b6/B0_55 ;
  wire  \inst_dob_mux_b6/B0_56 ;
  wire  \inst_dob_mux_b6/B0_57 ;
  wire  \inst_dob_mux_b6/B0_58 ;
  wire  \inst_dob_mux_b6/B0_59 ;
  wire  \inst_dob_mux_b6/B0_6 ;
  wire  \inst_dob_mux_b6/B0_60 ;
  wire  \inst_dob_mux_b6/B0_61 ;
  wire  \inst_dob_mux_b6/B0_62 ;
  wire  \inst_dob_mux_b6/B0_63 ;
  wire  \inst_dob_mux_b6/B0_7 ;
  wire  \inst_dob_mux_b6/B0_8 ;
  wire  \inst_dob_mux_b6/B0_9 ;
  wire  \inst_dob_mux_b6/B1_0 ;
  wire  \inst_dob_mux_b6/B1_1 ;
  wire  \inst_dob_mux_b6/B1_10 ;
  wire  \inst_dob_mux_b6/B1_11 ;
  wire  \inst_dob_mux_b6/B1_12 ;
  wire  \inst_dob_mux_b6/B1_13 ;
  wire  \inst_dob_mux_b6/B1_14 ;
  wire  \inst_dob_mux_b6/B1_15 ;
  wire  \inst_dob_mux_b6/B1_16 ;
  wire  \inst_dob_mux_b6/B1_17 ;
  wire  \inst_dob_mux_b6/B1_18 ;
  wire  \inst_dob_mux_b6/B1_19 ;
  wire  \inst_dob_mux_b6/B1_2 ;
  wire  \inst_dob_mux_b6/B1_20 ;
  wire  \inst_dob_mux_b6/B1_21 ;
  wire  \inst_dob_mux_b6/B1_22 ;
  wire  \inst_dob_mux_b6/B1_23 ;
  wire  \inst_dob_mux_b6/B1_24 ;
  wire  \inst_dob_mux_b6/B1_25 ;
  wire  \inst_dob_mux_b6/B1_26 ;
  wire  \inst_dob_mux_b6/B1_27 ;
  wire  \inst_dob_mux_b6/B1_28 ;
  wire  \inst_dob_mux_b6/B1_29 ;
  wire  \inst_dob_mux_b6/B1_3 ;
  wire  \inst_dob_mux_b6/B1_30 ;
  wire  \inst_dob_mux_b6/B1_31 ;
  wire  \inst_dob_mux_b6/B1_4 ;
  wire  \inst_dob_mux_b6/B1_5 ;
  wire  \inst_dob_mux_b6/B1_6 ;
  wire  \inst_dob_mux_b6/B1_7 ;
  wire  \inst_dob_mux_b6/B1_8 ;
  wire  \inst_dob_mux_b6/B1_9 ;
  wire  \inst_dob_mux_b6/B2_0 ;
  wire  \inst_dob_mux_b6/B2_1 ;
  wire  \inst_dob_mux_b6/B2_10 ;
  wire  \inst_dob_mux_b6/B2_11 ;
  wire  \inst_dob_mux_b6/B2_12 ;
  wire  \inst_dob_mux_b6/B2_13 ;
  wire  \inst_dob_mux_b6/B2_14 ;
  wire  \inst_dob_mux_b6/B2_15 ;
  wire  \inst_dob_mux_b6/B2_2 ;
  wire  \inst_dob_mux_b6/B2_3 ;
  wire  \inst_dob_mux_b6/B2_4 ;
  wire  \inst_dob_mux_b6/B2_5 ;
  wire  \inst_dob_mux_b6/B2_6 ;
  wire  \inst_dob_mux_b6/B2_7 ;
  wire  \inst_dob_mux_b6/B2_8 ;
  wire  \inst_dob_mux_b6/B2_9 ;
  wire  \inst_dob_mux_b6/B3_0 ;
  wire  \inst_dob_mux_b6/B3_1 ;
  wire  \inst_dob_mux_b6/B3_2 ;
  wire  \inst_dob_mux_b6/B3_3 ;
  wire  \inst_dob_mux_b6/B3_4 ;
  wire  \inst_dob_mux_b6/B3_5 ;
  wire  \inst_dob_mux_b6/B3_6 ;
  wire  \inst_dob_mux_b6/B3_7 ;
  wire  \inst_dob_mux_b6/B4_0 ;
  wire  \inst_dob_mux_b6/B4_1 ;
  wire  \inst_dob_mux_b6/B4_2 ;
  wire  \inst_dob_mux_b6/B4_3 ;
  wire  \inst_dob_mux_b6/B5_0 ;
  wire  \inst_dob_mux_b6/B5_1 ;
  wire  \inst_dob_mux_b7/B0_0 ;
  wire  \inst_dob_mux_b7/B0_1 ;
  wire  \inst_dob_mux_b7/B0_10 ;
  wire  \inst_dob_mux_b7/B0_11 ;
  wire  \inst_dob_mux_b7/B0_12 ;
  wire  \inst_dob_mux_b7/B0_13 ;
  wire  \inst_dob_mux_b7/B0_14 ;
  wire  \inst_dob_mux_b7/B0_15 ;
  wire  \inst_dob_mux_b7/B0_16 ;
  wire  \inst_dob_mux_b7/B0_17 ;
  wire  \inst_dob_mux_b7/B0_18 ;
  wire  \inst_dob_mux_b7/B0_19 ;
  wire  \inst_dob_mux_b7/B0_2 ;
  wire  \inst_dob_mux_b7/B0_20 ;
  wire  \inst_dob_mux_b7/B0_21 ;
  wire  \inst_dob_mux_b7/B0_22 ;
  wire  \inst_dob_mux_b7/B0_23 ;
  wire  \inst_dob_mux_b7/B0_24 ;
  wire  \inst_dob_mux_b7/B0_25 ;
  wire  \inst_dob_mux_b7/B0_26 ;
  wire  \inst_dob_mux_b7/B0_27 ;
  wire  \inst_dob_mux_b7/B0_28 ;
  wire  \inst_dob_mux_b7/B0_29 ;
  wire  \inst_dob_mux_b7/B0_3 ;
  wire  \inst_dob_mux_b7/B0_30 ;
  wire  \inst_dob_mux_b7/B0_31 ;
  wire  \inst_dob_mux_b7/B0_32 ;
  wire  \inst_dob_mux_b7/B0_33 ;
  wire  \inst_dob_mux_b7/B0_34 ;
  wire  \inst_dob_mux_b7/B0_35 ;
  wire  \inst_dob_mux_b7/B0_36 ;
  wire  \inst_dob_mux_b7/B0_37 ;
  wire  \inst_dob_mux_b7/B0_38 ;
  wire  \inst_dob_mux_b7/B0_39 ;
  wire  \inst_dob_mux_b7/B0_4 ;
  wire  \inst_dob_mux_b7/B0_40 ;
  wire  \inst_dob_mux_b7/B0_41 ;
  wire  \inst_dob_mux_b7/B0_42 ;
  wire  \inst_dob_mux_b7/B0_43 ;
  wire  \inst_dob_mux_b7/B0_44 ;
  wire  \inst_dob_mux_b7/B0_45 ;
  wire  \inst_dob_mux_b7/B0_46 ;
  wire  \inst_dob_mux_b7/B0_47 ;
  wire  \inst_dob_mux_b7/B0_48 ;
  wire  \inst_dob_mux_b7/B0_49 ;
  wire  \inst_dob_mux_b7/B0_5 ;
  wire  \inst_dob_mux_b7/B0_50 ;
  wire  \inst_dob_mux_b7/B0_51 ;
  wire  \inst_dob_mux_b7/B0_52 ;
  wire  \inst_dob_mux_b7/B0_53 ;
  wire  \inst_dob_mux_b7/B0_54 ;
  wire  \inst_dob_mux_b7/B0_55 ;
  wire  \inst_dob_mux_b7/B0_56 ;
  wire  \inst_dob_mux_b7/B0_57 ;
  wire  \inst_dob_mux_b7/B0_58 ;
  wire  \inst_dob_mux_b7/B0_59 ;
  wire  \inst_dob_mux_b7/B0_6 ;
  wire  \inst_dob_mux_b7/B0_60 ;
  wire  \inst_dob_mux_b7/B0_61 ;
  wire  \inst_dob_mux_b7/B0_62 ;
  wire  \inst_dob_mux_b7/B0_63 ;
  wire  \inst_dob_mux_b7/B0_7 ;
  wire  \inst_dob_mux_b7/B0_8 ;
  wire  \inst_dob_mux_b7/B0_9 ;
  wire  \inst_dob_mux_b7/B1_0 ;
  wire  \inst_dob_mux_b7/B1_1 ;
  wire  \inst_dob_mux_b7/B1_10 ;
  wire  \inst_dob_mux_b7/B1_11 ;
  wire  \inst_dob_mux_b7/B1_12 ;
  wire  \inst_dob_mux_b7/B1_13 ;
  wire  \inst_dob_mux_b7/B1_14 ;
  wire  \inst_dob_mux_b7/B1_15 ;
  wire  \inst_dob_mux_b7/B1_16 ;
  wire  \inst_dob_mux_b7/B1_17 ;
  wire  \inst_dob_mux_b7/B1_18 ;
  wire  \inst_dob_mux_b7/B1_19 ;
  wire  \inst_dob_mux_b7/B1_2 ;
  wire  \inst_dob_mux_b7/B1_20 ;
  wire  \inst_dob_mux_b7/B1_21 ;
  wire  \inst_dob_mux_b7/B1_22 ;
  wire  \inst_dob_mux_b7/B1_23 ;
  wire  \inst_dob_mux_b7/B1_24 ;
  wire  \inst_dob_mux_b7/B1_25 ;
  wire  \inst_dob_mux_b7/B1_26 ;
  wire  \inst_dob_mux_b7/B1_27 ;
  wire  \inst_dob_mux_b7/B1_28 ;
  wire  \inst_dob_mux_b7/B1_29 ;
  wire  \inst_dob_mux_b7/B1_3 ;
  wire  \inst_dob_mux_b7/B1_30 ;
  wire  \inst_dob_mux_b7/B1_31 ;
  wire  \inst_dob_mux_b7/B1_4 ;
  wire  \inst_dob_mux_b7/B1_5 ;
  wire  \inst_dob_mux_b7/B1_6 ;
  wire  \inst_dob_mux_b7/B1_7 ;
  wire  \inst_dob_mux_b7/B1_8 ;
  wire  \inst_dob_mux_b7/B1_9 ;
  wire  \inst_dob_mux_b7/B2_0 ;
  wire  \inst_dob_mux_b7/B2_1 ;
  wire  \inst_dob_mux_b7/B2_10 ;
  wire  \inst_dob_mux_b7/B2_11 ;
  wire  \inst_dob_mux_b7/B2_12 ;
  wire  \inst_dob_mux_b7/B2_13 ;
  wire  \inst_dob_mux_b7/B2_14 ;
  wire  \inst_dob_mux_b7/B2_15 ;
  wire  \inst_dob_mux_b7/B2_2 ;
  wire  \inst_dob_mux_b7/B2_3 ;
  wire  \inst_dob_mux_b7/B2_4 ;
  wire  \inst_dob_mux_b7/B2_5 ;
  wire  \inst_dob_mux_b7/B2_6 ;
  wire  \inst_dob_mux_b7/B2_7 ;
  wire  \inst_dob_mux_b7/B2_8 ;
  wire  \inst_dob_mux_b7/B2_9 ;
  wire  \inst_dob_mux_b7/B3_0 ;
  wire  \inst_dob_mux_b7/B3_1 ;
  wire  \inst_dob_mux_b7/B3_2 ;
  wire  \inst_dob_mux_b7/B3_3 ;
  wire  \inst_dob_mux_b7/B3_4 ;
  wire  \inst_dob_mux_b7/B3_5 ;
  wire  \inst_dob_mux_b7/B3_6 ;
  wire  \inst_dob_mux_b7/B3_7 ;
  wire  \inst_dob_mux_b7/B4_0 ;
  wire  \inst_dob_mux_b7/B4_1 ;
  wire  \inst_dob_mux_b7/B4_2 ;
  wire  \inst_dob_mux_b7/B4_3 ;
  wire  \inst_dob_mux_b7/B5_0 ;
  wire  \inst_dob_mux_b7/B5_1 ;
  wire  \inst_dob_mux_b8/B0_0 ;
  wire  \inst_dob_mux_b8/B0_1 ;
  wire  \inst_dob_mux_b8/B0_10 ;
  wire  \inst_dob_mux_b8/B0_11 ;
  wire  \inst_dob_mux_b8/B0_12 ;
  wire  \inst_dob_mux_b8/B0_13 ;
  wire  \inst_dob_mux_b8/B0_14 ;
  wire  \inst_dob_mux_b8/B0_15 ;
  wire  \inst_dob_mux_b8/B0_16 ;
  wire  \inst_dob_mux_b8/B0_17 ;
  wire  \inst_dob_mux_b8/B0_18 ;
  wire  \inst_dob_mux_b8/B0_19 ;
  wire  \inst_dob_mux_b8/B0_2 ;
  wire  \inst_dob_mux_b8/B0_20 ;
  wire  \inst_dob_mux_b8/B0_21 ;
  wire  \inst_dob_mux_b8/B0_22 ;
  wire  \inst_dob_mux_b8/B0_23 ;
  wire  \inst_dob_mux_b8/B0_24 ;
  wire  \inst_dob_mux_b8/B0_25 ;
  wire  \inst_dob_mux_b8/B0_26 ;
  wire  \inst_dob_mux_b8/B0_27 ;
  wire  \inst_dob_mux_b8/B0_28 ;
  wire  \inst_dob_mux_b8/B0_29 ;
  wire  \inst_dob_mux_b8/B0_3 ;
  wire  \inst_dob_mux_b8/B0_30 ;
  wire  \inst_dob_mux_b8/B0_31 ;
  wire  \inst_dob_mux_b8/B0_32 ;
  wire  \inst_dob_mux_b8/B0_33 ;
  wire  \inst_dob_mux_b8/B0_34 ;
  wire  \inst_dob_mux_b8/B0_35 ;
  wire  \inst_dob_mux_b8/B0_36 ;
  wire  \inst_dob_mux_b8/B0_37 ;
  wire  \inst_dob_mux_b8/B0_38 ;
  wire  \inst_dob_mux_b8/B0_39 ;
  wire  \inst_dob_mux_b8/B0_4 ;
  wire  \inst_dob_mux_b8/B0_40 ;
  wire  \inst_dob_mux_b8/B0_41 ;
  wire  \inst_dob_mux_b8/B0_42 ;
  wire  \inst_dob_mux_b8/B0_43 ;
  wire  \inst_dob_mux_b8/B0_44 ;
  wire  \inst_dob_mux_b8/B0_45 ;
  wire  \inst_dob_mux_b8/B0_46 ;
  wire  \inst_dob_mux_b8/B0_47 ;
  wire  \inst_dob_mux_b8/B0_48 ;
  wire  \inst_dob_mux_b8/B0_49 ;
  wire  \inst_dob_mux_b8/B0_5 ;
  wire  \inst_dob_mux_b8/B0_50 ;
  wire  \inst_dob_mux_b8/B0_51 ;
  wire  \inst_dob_mux_b8/B0_52 ;
  wire  \inst_dob_mux_b8/B0_53 ;
  wire  \inst_dob_mux_b8/B0_54 ;
  wire  \inst_dob_mux_b8/B0_55 ;
  wire  \inst_dob_mux_b8/B0_56 ;
  wire  \inst_dob_mux_b8/B0_57 ;
  wire  \inst_dob_mux_b8/B0_58 ;
  wire  \inst_dob_mux_b8/B0_59 ;
  wire  \inst_dob_mux_b8/B0_6 ;
  wire  \inst_dob_mux_b8/B0_60 ;
  wire  \inst_dob_mux_b8/B0_61 ;
  wire  \inst_dob_mux_b8/B0_62 ;
  wire  \inst_dob_mux_b8/B0_63 ;
  wire  \inst_dob_mux_b8/B0_7 ;
  wire  \inst_dob_mux_b8/B0_8 ;
  wire  \inst_dob_mux_b8/B0_9 ;
  wire  \inst_dob_mux_b8/B1_0 ;
  wire  \inst_dob_mux_b8/B1_1 ;
  wire  \inst_dob_mux_b8/B1_10 ;
  wire  \inst_dob_mux_b8/B1_11 ;
  wire  \inst_dob_mux_b8/B1_12 ;
  wire  \inst_dob_mux_b8/B1_13 ;
  wire  \inst_dob_mux_b8/B1_14 ;
  wire  \inst_dob_mux_b8/B1_15 ;
  wire  \inst_dob_mux_b8/B1_16 ;
  wire  \inst_dob_mux_b8/B1_17 ;
  wire  \inst_dob_mux_b8/B1_18 ;
  wire  \inst_dob_mux_b8/B1_19 ;
  wire  \inst_dob_mux_b8/B1_2 ;
  wire  \inst_dob_mux_b8/B1_20 ;
  wire  \inst_dob_mux_b8/B1_21 ;
  wire  \inst_dob_mux_b8/B1_22 ;
  wire  \inst_dob_mux_b8/B1_23 ;
  wire  \inst_dob_mux_b8/B1_24 ;
  wire  \inst_dob_mux_b8/B1_25 ;
  wire  \inst_dob_mux_b8/B1_26 ;
  wire  \inst_dob_mux_b8/B1_27 ;
  wire  \inst_dob_mux_b8/B1_28 ;
  wire  \inst_dob_mux_b8/B1_29 ;
  wire  \inst_dob_mux_b8/B1_3 ;
  wire  \inst_dob_mux_b8/B1_30 ;
  wire  \inst_dob_mux_b8/B1_31 ;
  wire  \inst_dob_mux_b8/B1_4 ;
  wire  \inst_dob_mux_b8/B1_5 ;
  wire  \inst_dob_mux_b8/B1_6 ;
  wire  \inst_dob_mux_b8/B1_7 ;
  wire  \inst_dob_mux_b8/B1_8 ;
  wire  \inst_dob_mux_b8/B1_9 ;
  wire  \inst_dob_mux_b8/B2_0 ;
  wire  \inst_dob_mux_b8/B2_1 ;
  wire  \inst_dob_mux_b8/B2_10 ;
  wire  \inst_dob_mux_b8/B2_11 ;
  wire  \inst_dob_mux_b8/B2_12 ;
  wire  \inst_dob_mux_b8/B2_13 ;
  wire  \inst_dob_mux_b8/B2_14 ;
  wire  \inst_dob_mux_b8/B2_15 ;
  wire  \inst_dob_mux_b8/B2_2 ;
  wire  \inst_dob_mux_b8/B2_3 ;
  wire  \inst_dob_mux_b8/B2_4 ;
  wire  \inst_dob_mux_b8/B2_5 ;
  wire  \inst_dob_mux_b8/B2_6 ;
  wire  \inst_dob_mux_b8/B2_7 ;
  wire  \inst_dob_mux_b8/B2_8 ;
  wire  \inst_dob_mux_b8/B2_9 ;
  wire  \inst_dob_mux_b8/B3_0 ;
  wire  \inst_dob_mux_b8/B3_1 ;
  wire  \inst_dob_mux_b8/B3_2 ;
  wire  \inst_dob_mux_b8/B3_3 ;
  wire  \inst_dob_mux_b8/B3_4 ;
  wire  \inst_dob_mux_b8/B3_5 ;
  wire  \inst_dob_mux_b8/B3_6 ;
  wire  \inst_dob_mux_b8/B3_7 ;
  wire  \inst_dob_mux_b8/B4_0 ;
  wire  \inst_dob_mux_b8/B4_1 ;
  wire  \inst_dob_mux_b8/B4_2 ;
  wire  \inst_dob_mux_b8/B4_3 ;
  wire  \inst_dob_mux_b8/B5_0 ;
  wire  \inst_dob_mux_b8/B5_1 ;
  wire  \inst_dob_mux_b9/B0_0 ;
  wire  \inst_dob_mux_b9/B0_1 ;
  wire  \inst_dob_mux_b9/B0_10 ;
  wire  \inst_dob_mux_b9/B0_11 ;
  wire  \inst_dob_mux_b9/B0_12 ;
  wire  \inst_dob_mux_b9/B0_13 ;
  wire  \inst_dob_mux_b9/B0_14 ;
  wire  \inst_dob_mux_b9/B0_15 ;
  wire  \inst_dob_mux_b9/B0_16 ;
  wire  \inst_dob_mux_b9/B0_17 ;
  wire  \inst_dob_mux_b9/B0_18 ;
  wire  \inst_dob_mux_b9/B0_19 ;
  wire  \inst_dob_mux_b9/B0_2 ;
  wire  \inst_dob_mux_b9/B0_20 ;
  wire  \inst_dob_mux_b9/B0_21 ;
  wire  \inst_dob_mux_b9/B0_22 ;
  wire  \inst_dob_mux_b9/B0_23 ;
  wire  \inst_dob_mux_b9/B0_24 ;
  wire  \inst_dob_mux_b9/B0_25 ;
  wire  \inst_dob_mux_b9/B0_26 ;
  wire  \inst_dob_mux_b9/B0_27 ;
  wire  \inst_dob_mux_b9/B0_28 ;
  wire  \inst_dob_mux_b9/B0_29 ;
  wire  \inst_dob_mux_b9/B0_3 ;
  wire  \inst_dob_mux_b9/B0_30 ;
  wire  \inst_dob_mux_b9/B0_31 ;
  wire  \inst_dob_mux_b9/B0_32 ;
  wire  \inst_dob_mux_b9/B0_33 ;
  wire  \inst_dob_mux_b9/B0_34 ;
  wire  \inst_dob_mux_b9/B0_35 ;
  wire  \inst_dob_mux_b9/B0_36 ;
  wire  \inst_dob_mux_b9/B0_37 ;
  wire  \inst_dob_mux_b9/B0_38 ;
  wire  \inst_dob_mux_b9/B0_39 ;
  wire  \inst_dob_mux_b9/B0_4 ;
  wire  \inst_dob_mux_b9/B0_40 ;
  wire  \inst_dob_mux_b9/B0_41 ;
  wire  \inst_dob_mux_b9/B0_42 ;
  wire  \inst_dob_mux_b9/B0_43 ;
  wire  \inst_dob_mux_b9/B0_44 ;
  wire  \inst_dob_mux_b9/B0_45 ;
  wire  \inst_dob_mux_b9/B0_46 ;
  wire  \inst_dob_mux_b9/B0_47 ;
  wire  \inst_dob_mux_b9/B0_48 ;
  wire  \inst_dob_mux_b9/B0_49 ;
  wire  \inst_dob_mux_b9/B0_5 ;
  wire  \inst_dob_mux_b9/B0_50 ;
  wire  \inst_dob_mux_b9/B0_51 ;
  wire  \inst_dob_mux_b9/B0_52 ;
  wire  \inst_dob_mux_b9/B0_53 ;
  wire  \inst_dob_mux_b9/B0_54 ;
  wire  \inst_dob_mux_b9/B0_55 ;
  wire  \inst_dob_mux_b9/B0_56 ;
  wire  \inst_dob_mux_b9/B0_57 ;
  wire  \inst_dob_mux_b9/B0_58 ;
  wire  \inst_dob_mux_b9/B0_59 ;
  wire  \inst_dob_mux_b9/B0_6 ;
  wire  \inst_dob_mux_b9/B0_60 ;
  wire  \inst_dob_mux_b9/B0_61 ;
  wire  \inst_dob_mux_b9/B0_62 ;
  wire  \inst_dob_mux_b9/B0_63 ;
  wire  \inst_dob_mux_b9/B0_7 ;
  wire  \inst_dob_mux_b9/B0_8 ;
  wire  \inst_dob_mux_b9/B0_9 ;
  wire  \inst_dob_mux_b9/B1_0 ;
  wire  \inst_dob_mux_b9/B1_1 ;
  wire  \inst_dob_mux_b9/B1_10 ;
  wire  \inst_dob_mux_b9/B1_11 ;
  wire  \inst_dob_mux_b9/B1_12 ;
  wire  \inst_dob_mux_b9/B1_13 ;
  wire  \inst_dob_mux_b9/B1_14 ;
  wire  \inst_dob_mux_b9/B1_15 ;
  wire  \inst_dob_mux_b9/B1_16 ;
  wire  \inst_dob_mux_b9/B1_17 ;
  wire  \inst_dob_mux_b9/B1_18 ;
  wire  \inst_dob_mux_b9/B1_19 ;
  wire  \inst_dob_mux_b9/B1_2 ;
  wire  \inst_dob_mux_b9/B1_20 ;
  wire  \inst_dob_mux_b9/B1_21 ;
  wire  \inst_dob_mux_b9/B1_22 ;
  wire  \inst_dob_mux_b9/B1_23 ;
  wire  \inst_dob_mux_b9/B1_24 ;
  wire  \inst_dob_mux_b9/B1_25 ;
  wire  \inst_dob_mux_b9/B1_26 ;
  wire  \inst_dob_mux_b9/B1_27 ;
  wire  \inst_dob_mux_b9/B1_28 ;
  wire  \inst_dob_mux_b9/B1_29 ;
  wire  \inst_dob_mux_b9/B1_3 ;
  wire  \inst_dob_mux_b9/B1_30 ;
  wire  \inst_dob_mux_b9/B1_31 ;
  wire  \inst_dob_mux_b9/B1_4 ;
  wire  \inst_dob_mux_b9/B1_5 ;
  wire  \inst_dob_mux_b9/B1_6 ;
  wire  \inst_dob_mux_b9/B1_7 ;
  wire  \inst_dob_mux_b9/B1_8 ;
  wire  \inst_dob_mux_b9/B1_9 ;
  wire  \inst_dob_mux_b9/B2_0 ;
  wire  \inst_dob_mux_b9/B2_1 ;
  wire  \inst_dob_mux_b9/B2_10 ;
  wire  \inst_dob_mux_b9/B2_11 ;
  wire  \inst_dob_mux_b9/B2_12 ;
  wire  \inst_dob_mux_b9/B2_13 ;
  wire  \inst_dob_mux_b9/B2_14 ;
  wire  \inst_dob_mux_b9/B2_15 ;
  wire  \inst_dob_mux_b9/B2_2 ;
  wire  \inst_dob_mux_b9/B2_3 ;
  wire  \inst_dob_mux_b9/B2_4 ;
  wire  \inst_dob_mux_b9/B2_5 ;
  wire  \inst_dob_mux_b9/B2_6 ;
  wire  \inst_dob_mux_b9/B2_7 ;
  wire  \inst_dob_mux_b9/B2_8 ;
  wire  \inst_dob_mux_b9/B2_9 ;
  wire  \inst_dob_mux_b9/B3_0 ;
  wire  \inst_dob_mux_b9/B3_1 ;
  wire  \inst_dob_mux_b9/B3_2 ;
  wire  \inst_dob_mux_b9/B3_3 ;
  wire  \inst_dob_mux_b9/B3_4 ;
  wire  \inst_dob_mux_b9/B3_5 ;
  wire  \inst_dob_mux_b9/B3_6 ;
  wire  \inst_dob_mux_b9/B3_7 ;
  wire  \inst_dob_mux_b9/B4_0 ;
  wire  \inst_dob_mux_b9/B4_1 ;
  wire  \inst_dob_mux_b9/B4_2 ;
  wire  \inst_dob_mux_b9/B4_3 ;
  wire  \inst_dob_mux_b9/B5_0 ;
  wire  \inst_dob_mux_b9/B5_1 ;
  wire and_Naddra$11$_Naddr_o;
  wire and_Naddra$11$_Naddr_o_and_cea;
  wire and_Naddra$12$_Naddr_o;
  wire and_Naddra$12$_Naddr_o_al_n54;
  wire and_Naddra$12$_addra_o;
  wire and_Naddra$12$_addra_o_al_n86;
  wire and_Naddrb$11$_Naddr_o;
  wire and_Naddrb$11$_Naddr_o_and_ceb;
  wire and_Naddrb$12$_Naddr_o;
  wire and_Naddrb$12$_Naddr_o_al_n57;
  wire and_Naddrb$12$_addrb_o;
  wire and_Naddrb$12$_addrb_o_al_n89;
  wire and_addra$12$_Naddra_o;
  wire and_addra$12$_Naddra_o_al_n70;
  wire and_addra$12$_addra$_o;
  wire and_addra$12$_addra$_o_al_n102;
  wire and_addrb$12$_Naddrb_o;
  wire and_addrb$12$_Naddrb_o_al_n73;
  wire and_addrb$12$_addrb$_o;
  wire and_addrb$12$_addrb$_o_al_n105;
  wire inst_dob_i0_000;
  wire inst_dob_i0_001;
  wire inst_dob_i0_002;
  wire inst_dob_i0_003;
  wire inst_dob_i0_004;
  wire inst_dob_i0_005;
  wire inst_dob_i0_006;
  wire inst_dob_i0_007;
  wire inst_dob_i0_008;
  wire inst_dob_i0_009;
  wire inst_dob_i0_010;
  wire inst_dob_i0_011;
  wire inst_dob_i0_012;
  wire inst_dob_i0_013;
  wire inst_dob_i0_014;
  wire inst_dob_i0_015;
  wire inst_dob_i10_000;
  wire inst_dob_i10_001;
  wire inst_dob_i10_002;
  wire inst_dob_i10_003;
  wire inst_dob_i10_004;
  wire inst_dob_i10_005;
  wire inst_dob_i10_006;
  wire inst_dob_i10_007;
  wire inst_dob_i10_008;
  wire inst_dob_i12_000;
  wire inst_dob_i12_001;
  wire inst_dob_i12_002;
  wire inst_dob_i12_003;
  wire inst_dob_i12_004;
  wire inst_dob_i12_005;
  wire inst_dob_i12_006;
  wire inst_dob_i12_007;
  wire inst_dob_i12_008;
  wire inst_dob_i14_000;
  wire inst_dob_i14_001;
  wire inst_dob_i14_002;
  wire inst_dob_i14_003;
  wire inst_dob_i14_004;
  wire inst_dob_i14_005;
  wire inst_dob_i14_006;
  wire inst_dob_i14_007;
  wire inst_dob_i14_008;
  wire inst_dob_i16_000;
  wire inst_dob_i16_001;
  wire inst_dob_i16_002;
  wire inst_dob_i16_003;
  wire inst_dob_i16_004;
  wire inst_dob_i16_005;
  wire inst_dob_i16_006;
  wire inst_dob_i16_007;
  wire inst_dob_i16_008;
  wire inst_dob_i16_009;
  wire inst_dob_i16_010;
  wire inst_dob_i16_011;
  wire inst_dob_i16_012;
  wire inst_dob_i16_013;
  wire inst_dob_i16_014;
  wire inst_dob_i16_015;
  wire inst_dob_i18_000;
  wire inst_dob_i18_001;
  wire inst_dob_i18_002;
  wire inst_dob_i18_003;
  wire inst_dob_i18_004;
  wire inst_dob_i18_005;
  wire inst_dob_i18_006;
  wire inst_dob_i18_007;
  wire inst_dob_i18_008;
  wire inst_dob_i20_000;
  wire inst_dob_i20_001;
  wire inst_dob_i20_002;
  wire inst_dob_i20_003;
  wire inst_dob_i20_004;
  wire inst_dob_i20_005;
  wire inst_dob_i20_006;
  wire inst_dob_i20_007;
  wire inst_dob_i20_008;
  wire inst_dob_i22_000;
  wire inst_dob_i22_001;
  wire inst_dob_i22_002;
  wire inst_dob_i22_003;
  wire inst_dob_i22_004;
  wire inst_dob_i22_005;
  wire inst_dob_i22_006;
  wire inst_dob_i22_007;
  wire inst_dob_i22_008;
  wire inst_dob_i24_000;
  wire inst_dob_i24_001;
  wire inst_dob_i24_002;
  wire inst_dob_i24_003;
  wire inst_dob_i24_004;
  wire inst_dob_i24_005;
  wire inst_dob_i24_006;
  wire inst_dob_i24_007;
  wire inst_dob_i24_008;
  wire inst_dob_i26_000;
  wire inst_dob_i26_001;
  wire inst_dob_i26_002;
  wire inst_dob_i26_003;
  wire inst_dob_i26_004;
  wire inst_dob_i26_005;
  wire inst_dob_i26_006;
  wire inst_dob_i26_007;
  wire inst_dob_i26_008;
  wire inst_dob_i28_000;
  wire inst_dob_i28_001;
  wire inst_dob_i28_002;
  wire inst_dob_i28_003;
  wire inst_dob_i28_004;
  wire inst_dob_i28_005;
  wire inst_dob_i28_006;
  wire inst_dob_i28_007;
  wire inst_dob_i28_008;
  wire inst_dob_i2_000;
  wire inst_dob_i2_001;
  wire inst_dob_i2_002;
  wire inst_dob_i2_003;
  wire inst_dob_i2_004;
  wire inst_dob_i2_005;
  wire inst_dob_i2_006;
  wire inst_dob_i2_007;
  wire inst_dob_i2_008;
  wire inst_dob_i30_000;
  wire inst_dob_i30_001;
  wire inst_dob_i30_002;
  wire inst_dob_i30_003;
  wire inst_dob_i30_004;
  wire inst_dob_i30_005;
  wire inst_dob_i30_006;
  wire inst_dob_i30_007;
  wire inst_dob_i30_008;
  wire inst_dob_i32_000;
  wire inst_dob_i32_001;
  wire inst_dob_i32_002;
  wire inst_dob_i32_003;
  wire inst_dob_i32_004;
  wire inst_dob_i32_005;
  wire inst_dob_i32_006;
  wire inst_dob_i32_007;
  wire inst_dob_i32_008;
  wire inst_dob_i32_009;
  wire inst_dob_i32_010;
  wire inst_dob_i32_011;
  wire inst_dob_i32_012;
  wire inst_dob_i32_013;
  wire inst_dob_i32_014;
  wire inst_dob_i32_015;
  wire inst_dob_i34_000;
  wire inst_dob_i34_001;
  wire inst_dob_i34_002;
  wire inst_dob_i34_003;
  wire inst_dob_i34_004;
  wire inst_dob_i34_005;
  wire inst_dob_i34_006;
  wire inst_dob_i34_007;
  wire inst_dob_i34_008;
  wire inst_dob_i36_000;
  wire inst_dob_i36_001;
  wire inst_dob_i36_002;
  wire inst_dob_i36_003;
  wire inst_dob_i36_004;
  wire inst_dob_i36_005;
  wire inst_dob_i36_006;
  wire inst_dob_i36_007;
  wire inst_dob_i36_008;
  wire inst_dob_i38_000;
  wire inst_dob_i38_001;
  wire inst_dob_i38_002;
  wire inst_dob_i38_003;
  wire inst_dob_i38_004;
  wire inst_dob_i38_005;
  wire inst_dob_i38_006;
  wire inst_dob_i38_007;
  wire inst_dob_i38_008;
  wire inst_dob_i40_000;
  wire inst_dob_i40_001;
  wire inst_dob_i40_002;
  wire inst_dob_i40_003;
  wire inst_dob_i40_004;
  wire inst_dob_i40_005;
  wire inst_dob_i40_006;
  wire inst_dob_i40_007;
  wire inst_dob_i40_008;
  wire inst_dob_i42_000;
  wire inst_dob_i42_001;
  wire inst_dob_i42_002;
  wire inst_dob_i42_003;
  wire inst_dob_i42_004;
  wire inst_dob_i42_005;
  wire inst_dob_i42_006;
  wire inst_dob_i42_007;
  wire inst_dob_i42_008;
  wire inst_dob_i44_000;
  wire inst_dob_i44_001;
  wire inst_dob_i44_002;
  wire inst_dob_i44_003;
  wire inst_dob_i44_004;
  wire inst_dob_i44_005;
  wire inst_dob_i44_006;
  wire inst_dob_i44_007;
  wire inst_dob_i44_008;
  wire inst_dob_i46_000;
  wire inst_dob_i46_001;
  wire inst_dob_i46_002;
  wire inst_dob_i46_003;
  wire inst_dob_i46_004;
  wire inst_dob_i46_005;
  wire inst_dob_i46_006;
  wire inst_dob_i46_007;
  wire inst_dob_i46_008;
  wire inst_dob_i48_000;
  wire inst_dob_i48_001;
  wire inst_dob_i48_002;
  wire inst_dob_i48_003;
  wire inst_dob_i48_004;
  wire inst_dob_i48_005;
  wire inst_dob_i48_006;
  wire inst_dob_i48_007;
  wire inst_dob_i48_008;
  wire inst_dob_i48_009;
  wire inst_dob_i48_010;
  wire inst_dob_i48_011;
  wire inst_dob_i48_012;
  wire inst_dob_i48_013;
  wire inst_dob_i48_014;
  wire inst_dob_i48_015;
  wire inst_dob_i4_000;
  wire inst_dob_i4_001;
  wire inst_dob_i4_002;
  wire inst_dob_i4_003;
  wire inst_dob_i4_004;
  wire inst_dob_i4_005;
  wire inst_dob_i4_006;
  wire inst_dob_i4_007;
  wire inst_dob_i4_008;
  wire inst_dob_i50_000;
  wire inst_dob_i50_001;
  wire inst_dob_i50_002;
  wire inst_dob_i50_003;
  wire inst_dob_i50_004;
  wire inst_dob_i50_005;
  wire inst_dob_i50_006;
  wire inst_dob_i50_007;
  wire inst_dob_i50_008;
  wire inst_dob_i52_000;
  wire inst_dob_i52_001;
  wire inst_dob_i52_002;
  wire inst_dob_i52_003;
  wire inst_dob_i52_004;
  wire inst_dob_i52_005;
  wire inst_dob_i52_006;
  wire inst_dob_i52_007;
  wire inst_dob_i52_008;
  wire inst_dob_i54_000;
  wire inst_dob_i54_001;
  wire inst_dob_i54_002;
  wire inst_dob_i54_003;
  wire inst_dob_i54_004;
  wire inst_dob_i54_005;
  wire inst_dob_i54_006;
  wire inst_dob_i54_007;
  wire inst_dob_i54_008;
  wire inst_dob_i56_000;
  wire inst_dob_i56_001;
  wire inst_dob_i56_002;
  wire inst_dob_i56_003;
  wire inst_dob_i56_004;
  wire inst_dob_i56_005;
  wire inst_dob_i56_006;
  wire inst_dob_i56_007;
  wire inst_dob_i56_008;
  wire inst_dob_i58_000;
  wire inst_dob_i58_001;
  wire inst_dob_i58_002;
  wire inst_dob_i58_003;
  wire inst_dob_i58_004;
  wire inst_dob_i58_005;
  wire inst_dob_i58_006;
  wire inst_dob_i58_007;
  wire inst_dob_i58_008;
  wire inst_dob_i60_000;
  wire inst_dob_i60_001;
  wire inst_dob_i60_002;
  wire inst_dob_i60_003;
  wire inst_dob_i60_004;
  wire inst_dob_i60_005;
  wire inst_dob_i60_006;
  wire inst_dob_i60_007;
  wire inst_dob_i60_008;
  wire inst_dob_i62_000;
  wire inst_dob_i62_001;
  wire inst_dob_i62_002;
  wire inst_dob_i62_003;
  wire inst_dob_i62_004;
  wire inst_dob_i62_005;
  wire inst_dob_i62_006;
  wire inst_dob_i62_007;
  wire inst_dob_i62_008;
  wire inst_dob_i64_000;
  wire inst_dob_i64_001;
  wire inst_dob_i64_002;
  wire inst_dob_i64_003;
  wire inst_dob_i64_004;
  wire inst_dob_i64_005;
  wire inst_dob_i64_006;
  wire inst_dob_i64_007;
  wire inst_dob_i64_008;
  wire inst_dob_i64_009;
  wire inst_dob_i64_010;
  wire inst_dob_i64_011;
  wire inst_dob_i64_012;
  wire inst_dob_i64_013;
  wire inst_dob_i64_014;
  wire inst_dob_i64_015;
  wire inst_dob_i6_000;
  wire inst_dob_i6_001;
  wire inst_dob_i6_002;
  wire inst_dob_i6_003;
  wire inst_dob_i6_004;
  wire inst_dob_i6_005;
  wire inst_dob_i6_006;
  wire inst_dob_i6_007;
  wire inst_dob_i6_008;
  wire inst_dob_i8_000;
  wire inst_dob_i8_001;
  wire inst_dob_i8_002;
  wire inst_dob_i8_003;
  wire inst_dob_i8_004;
  wire inst_dob_i8_005;
  wire inst_dob_i8_006;
  wire inst_dob_i8_007;
  wire inst_dob_i8_008;

  reg_sr_as_w1 addrb_pipe_b0 (
    .clk(clkb),
    .d(addrb[9]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[0]));
  reg_sr_as_w1 addrb_pipe_b1 (
    .clk(clkb),
    .d(addrb[10]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[1]));
  reg_sr_as_w1 addrb_pipe_b2 (
    .clk(clkb),
    .d(addrb[11]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[2]));
  reg_sr_as_w1 addrb_pipe_b3 (
    .clk(clkb),
    .d(addrb[12]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[3]));
  reg_sr_as_w1 addrb_pipe_b4 (
    .clk(clkb),
    .d(addrb[13]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[4]));
  reg_sr_as_w1 addrb_pipe_b5 (
    .clk(clkb),
    .d(addrb[14]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[5]));
  reg_sr_as_w1 addrb_pipe_b6 (
    .clk(clkb),
    .d(addrb[15]),
    .en(ceb),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped[6]));
  and and_Naddra$11$_Naddr_o_and_cea_i (and_Naddra$11$_Naddr_o_and_cea, and_Naddra$11$_Naddr_o, cea);
  and \and_Naddra[11]_Naddr  (and_Naddra$11$_Naddr_o, ~addra[11], ~addra[12], ~addra[13], ~addra[14], addra[15]);
  and \and_Naddra[12]_Naddr  (and_Naddra$12$_Naddr_o, ~addra[12], ~addra[13], ~addra[14], ~addra[15]);
  and \and_Naddra[12]_Naddr_al_u54  (and_Naddra$12$_Naddr_o_al_n54, ~addra[12], ~addra[13], addra[14], ~addra[15]);
  and \and_Naddra[12]_addra  (and_Naddra$12$_addra_o, ~addra[12], addra[13], ~addra[14], ~addra[15]);
  and \and_Naddra[12]_addra_al_u86  (and_Naddra$12$_addra_o_al_n86, ~addra[12], addra[13], addra[14], ~addra[15]);
  and and_Naddrb$11$_Naddr_o_and_ceb_i (and_Naddrb$11$_Naddr_o_and_ceb, and_Naddrb$11$_Naddr_o, ceb);
  and \and_Naddrb[11]_Naddr  (and_Naddrb$11$_Naddr_o, ~addrb[11], ~addrb[12], ~addrb[13], ~addrb[14], addrb[15]);
  and \and_Naddrb[12]_Naddr  (and_Naddrb$12$_Naddr_o, ~addrb[12], ~addrb[13], ~addrb[14], ~addrb[15]);
  and \and_Naddrb[12]_Naddr_al_u57  (and_Naddrb$12$_Naddr_o_al_n57, ~addrb[12], ~addrb[13], addrb[14], ~addrb[15]);
  and \and_Naddrb[12]_addrb  (and_Naddrb$12$_addrb_o, ~addrb[12], addrb[13], ~addrb[14], ~addrb[15]);
  and \and_Naddrb[12]_addrb_al_u89  (and_Naddrb$12$_addrb_o_al_n89, ~addrb[12], addrb[13], addrb[14], ~addrb[15]);
  and \and_addra[12]_Naddra  (and_addra$12$_Naddra_o, addra[12], ~addra[13], ~addra[14], ~addra[15]);
  and \and_addra[12]_Naddra_al_u70  (and_addra$12$_Naddra_o_al_n70, addra[12], ~addra[13], addra[14], ~addra[15]);
  and \and_addra[12]_addra[  (and_addra$12$_addra$_o, addra[12], addra[13], ~addra[14], ~addra[15]);
  and \and_addra[12]_addra[_al_u102  (and_addra$12$_addra$_o_al_n102, addra[12], addra[13], addra[14], ~addra[15]);
  and \and_addrb[12]_Naddrb  (and_addrb$12$_Naddrb_o, addrb[12], ~addrb[13], ~addrb[14], ~addrb[15]);
  and \and_addrb[12]_Naddrb_al_u73  (and_addrb$12$_Naddrb_o_al_n73, addrb[12], ~addrb[13], addrb[14], ~addrb[15]);
  and \and_addrb[12]_addrb[  (and_addrb$12$_addrb$_o, addrb[12], addrb[13], ~addrb[14], ~addrb[15]);
  and \and_addrb[12]_addrb[_al_u105  (and_addrb$12$_addrb$_o_al_n105, addrb[12], addrb[13], addrb[14], ~addrb[15]);
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_Naddr_o,addra[11:10]}),
    .csb({and_Naddrb$12$_Naddr_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i0_008,inst_dob_i0_007,inst_dob_i0_006,inst_dob_i0_005,inst_dob_i0_004,inst_dob_i0_003,inst_dob_i0_002,inst_dob_i0_001,inst_dob_i0_000}));
  // address_offset=0;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_009 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n69,open_n70,open_n71,open_n72,open_n73,open_n74,open_n75,dia[9],open_n76}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n99,open_n100,open_n101,open_n102,open_n103,open_n104,open_n105,open_n106,inst_dob_i0_009}));
  // address_offset=0;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_010 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n107,open_n108,open_n109,open_n110,open_n111,open_n112,open_n113,dia[10],open_n114}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n137,open_n138,open_n139,open_n140,open_n141,open_n142,open_n143,open_n144,inst_dob_i0_010}));
  // address_offset=0;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_011 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n145,open_n146,open_n147,open_n148,open_n149,open_n150,open_n151,dia[11],open_n152}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n175,open_n176,open_n177,open_n178,open_n179,open_n180,open_n181,open_n182,inst_dob_i0_011}));
  // address_offset=0;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_012 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n183,open_n184,open_n185,open_n186,open_n187,open_n188,open_n189,dia[12],open_n190}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n213,open_n214,open_n215,open_n216,open_n217,open_n218,open_n219,open_n220,inst_dob_i0_012}));
  // address_offset=0;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_013 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n221,open_n222,open_n223,open_n224,open_n225,open_n226,open_n227,dia[13],open_n228}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n251,open_n252,open_n253,open_n254,open_n255,open_n256,open_n257,open_n258,inst_dob_i0_013}));
  // address_offset=0;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_014 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n259,open_n260,open_n261,open_n262,open_n263,open_n264,open_n265,dia[14],open_n266}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n289,open_n290,open_n291,open_n292,open_n293,open_n294,open_n295,open_n296,inst_dob_i0_014}));
  // address_offset=0;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_015 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n297,open_n298,open_n299,open_n300,open_n301,open_n302,open_n303,dia[15],open_n304}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n327,open_n328,open_n329,open_n330,open_n331,open_n332,open_n333,open_n334,inst_dob_i0_015}));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_001024_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_Naddr_o,addra[11:10]}),
    .csb({and_Naddrb$12$_Naddr_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i2_008,inst_dob_i2_007,inst_dob_i2_006,inst_dob_i2_005,inst_dob_i2_004,inst_dob_i2_003,inst_dob_i2_002,inst_dob_i2_001,inst_dob_i2_000}));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_002048_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_Naddr_o,addra[11:10]}),
    .csb({and_Naddrb$12$_Naddr_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i4_008,inst_dob_i4_007,inst_dob_i4_006,inst_dob_i4_005,inst_dob_i4_004,inst_dob_i4_003,inst_dob_i4_002,inst_dob_i4_001,inst_dob_i4_000}));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_003072_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_Naddr_o,addra[11:10]}),
    .csb({and_Naddrb$12$_Naddr_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i6_008,inst_dob_i6_007,inst_dob_i6_006,inst_dob_i6_005,inst_dob_i6_004,inst_dob_i6_003,inst_dob_i6_002,inst_dob_i6_001,inst_dob_i6_000}));
  // address_offset=4096;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_004096_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_Naddra_o,addra[11:10]}),
    .csb({and_addrb$12$_Naddrb_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i8_008,inst_dob_i8_007,inst_dob_i8_006,inst_dob_i8_005,inst_dob_i8_004,inst_dob_i8_003,inst_dob_i8_002,inst_dob_i8_001,inst_dob_i8_000}));
  // address_offset=5120;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_005120_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_Naddra_o,addra[11:10]}),
    .csb({and_addrb$12$_Naddrb_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i10_008,inst_dob_i10_007,inst_dob_i10_006,inst_dob_i10_005,inst_dob_i10_004,inst_dob_i10_003,inst_dob_i10_002,inst_dob_i10_001,inst_dob_i10_000}));
  // address_offset=6144;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_006144_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_Naddra_o,addra[11:10]}),
    .csb({and_addrb$12$_Naddrb_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i12_008,inst_dob_i12_007,inst_dob_i12_006,inst_dob_i12_005,inst_dob_i12_004,inst_dob_i12_003,inst_dob_i12_002,inst_dob_i12_001,inst_dob_i12_000}));
  // address_offset=7168;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_007168_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_Naddra_o,addra[11:10]}),
    .csb({and_addrb$12$_Naddrb_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i14_008,inst_dob_i14_007,inst_dob_i14_006,inst_dob_i14_005,inst_dob_i14_004,inst_dob_i14_003,inst_dob_i14_002,inst_dob_i14_001,inst_dob_i14_000}));
  // address_offset=8192;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_addra_o,addra[11:10]}),
    .csb({and_Naddrb$12$_addrb_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i16_008,inst_dob_i16_007,inst_dob_i16_006,inst_dob_i16_005,inst_dob_i16_004,inst_dob_i16_003,inst_dob_i16_002,inst_dob_i16_001,inst_dob_i16_000}));
  // address_offset=8192;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_009 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n511,open_n512,open_n513,open_n514,open_n515,open_n516,open_n517,dia[9],open_n518}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n541,open_n542,open_n543,open_n544,open_n545,open_n546,open_n547,open_n548,inst_dob_i16_009}));
  // address_offset=8192;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_010 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n549,open_n550,open_n551,open_n552,open_n553,open_n554,open_n555,dia[10],open_n556}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n579,open_n580,open_n581,open_n582,open_n583,open_n584,open_n585,open_n586,inst_dob_i16_010}));
  // address_offset=8192;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_011 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n587,open_n588,open_n589,open_n590,open_n591,open_n592,open_n593,dia[11],open_n594}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n617,open_n618,open_n619,open_n620,open_n621,open_n622,open_n623,open_n624,inst_dob_i16_011}));
  // address_offset=8192;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_012 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n625,open_n626,open_n627,open_n628,open_n629,open_n630,open_n631,dia[12],open_n632}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n655,open_n656,open_n657,open_n658,open_n659,open_n660,open_n661,open_n662,inst_dob_i16_012}));
  // address_offset=8192;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_013 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n663,open_n664,open_n665,open_n666,open_n667,open_n668,open_n669,dia[13],open_n670}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n693,open_n694,open_n695,open_n696,open_n697,open_n698,open_n699,open_n700,inst_dob_i16_013}));
  // address_offset=8192;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_014 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n701,open_n702,open_n703,open_n704,open_n705,open_n706,open_n707,dia[14],open_n708}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n731,open_n732,open_n733,open_n734,open_n735,open_n736,open_n737,open_n738,inst_dob_i16_014}));
  // address_offset=8192;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_015 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n739,open_n740,open_n741,open_n742,open_n743,open_n744,open_n745,dia[15],open_n746}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n769,open_n770,open_n771,open_n772,open_n773,open_n774,open_n775,open_n776,inst_dob_i16_015}));
  // address_offset=9216;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_009216_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_addra_o,addra[11:10]}),
    .csb({and_Naddrb$12$_addrb_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i18_008,inst_dob_i18_007,inst_dob_i18_006,inst_dob_i18_005,inst_dob_i18_004,inst_dob_i18_003,inst_dob_i18_002,inst_dob_i18_001,inst_dob_i18_000}));
  // address_offset=10240;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_010240_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_addra_o,addra[11:10]}),
    .csb({and_Naddrb$12$_addrb_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i20_008,inst_dob_i20_007,inst_dob_i20_006,inst_dob_i20_005,inst_dob_i20_004,inst_dob_i20_003,inst_dob_i20_002,inst_dob_i20_001,inst_dob_i20_000}));
  // address_offset=11264;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_011264_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_addra_o,addra[11:10]}),
    .csb({and_Naddrb$12$_addrb_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i22_008,inst_dob_i22_007,inst_dob_i22_006,inst_dob_i22_005,inst_dob_i22_004,inst_dob_i22_003,inst_dob_i22_002,inst_dob_i22_001,inst_dob_i22_000}));
  // address_offset=12288;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_012288_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_addra$_o,addra[11:10]}),
    .csb({and_addrb$12$_addrb$_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i24_008,inst_dob_i24_007,inst_dob_i24_006,inst_dob_i24_005,inst_dob_i24_004,inst_dob_i24_003,inst_dob_i24_002,inst_dob_i24_001,inst_dob_i24_000}));
  // address_offset=13312;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_013312_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_addra$_o,addra[11:10]}),
    .csb({and_addrb$12$_addrb$_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i26_008,inst_dob_i26_007,inst_dob_i26_006,inst_dob_i26_005,inst_dob_i26_004,inst_dob_i26_003,inst_dob_i26_002,inst_dob_i26_001,inst_dob_i26_000}));
  // address_offset=14336;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_014336_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_addra$_o,addra[11:10]}),
    .csb({and_addrb$12$_addrb$_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i28_008,inst_dob_i28_007,inst_dob_i28_006,inst_dob_i28_005,inst_dob_i28_004,inst_dob_i28_003,inst_dob_i28_002,inst_dob_i28_001,inst_dob_i28_000}));
  // address_offset=15360;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_015360_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_addra$_o,addra[11:10]}),
    .csb({and_addrb$12$_addrb$_o,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i30_008,inst_dob_i30_007,inst_dob_i30_006,inst_dob_i30_005,inst_dob_i30_004,inst_dob_i30_003,inst_dob_i30_002,inst_dob_i30_001,inst_dob_i30_000}));
  // address_offset=16384;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_Naddr_o_al_n54,addra[11:10]}),
    .csb({and_Naddrb$12$_Naddr_o_al_n57,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i32_008,inst_dob_i32_007,inst_dob_i32_006,inst_dob_i32_005,inst_dob_i32_004,inst_dob_i32_003,inst_dob_i32_002,inst_dob_i32_001,inst_dob_i32_000}));
  // address_offset=16384;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_009 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n953,open_n954,open_n955,open_n956,open_n957,open_n958,open_n959,dia[9],open_n960}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n983,open_n984,open_n985,open_n986,open_n987,open_n988,open_n989,open_n990,inst_dob_i32_009}));
  // address_offset=16384;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_010 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n991,open_n992,open_n993,open_n994,open_n995,open_n996,open_n997,dia[10],open_n998}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1021,open_n1022,open_n1023,open_n1024,open_n1025,open_n1026,open_n1027,open_n1028,inst_dob_i32_010}));
  // address_offset=16384;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_011 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1029,open_n1030,open_n1031,open_n1032,open_n1033,open_n1034,open_n1035,dia[11],open_n1036}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1059,open_n1060,open_n1061,open_n1062,open_n1063,open_n1064,open_n1065,open_n1066,inst_dob_i32_011}));
  // address_offset=16384;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_012 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1067,open_n1068,open_n1069,open_n1070,open_n1071,open_n1072,open_n1073,dia[12],open_n1074}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1097,open_n1098,open_n1099,open_n1100,open_n1101,open_n1102,open_n1103,open_n1104,inst_dob_i32_012}));
  // address_offset=16384;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_013 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1105,open_n1106,open_n1107,open_n1108,open_n1109,open_n1110,open_n1111,dia[13],open_n1112}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1135,open_n1136,open_n1137,open_n1138,open_n1139,open_n1140,open_n1141,open_n1142,inst_dob_i32_013}));
  // address_offset=16384;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_014 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1143,open_n1144,open_n1145,open_n1146,open_n1147,open_n1148,open_n1149,dia[14],open_n1150}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1173,open_n1174,open_n1175,open_n1176,open_n1177,open_n1178,open_n1179,open_n1180,inst_dob_i32_014}));
  // address_offset=16384;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_015 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1181,open_n1182,open_n1183,open_n1184,open_n1185,open_n1186,open_n1187,dia[15],open_n1188}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1211,open_n1212,open_n1213,open_n1214,open_n1215,open_n1216,open_n1217,open_n1218,inst_dob_i32_015}));
  // address_offset=17408;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_017408_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_Naddr_o_al_n54,addra[11:10]}),
    .csb({and_Naddrb$12$_Naddr_o_al_n57,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i34_008,inst_dob_i34_007,inst_dob_i34_006,inst_dob_i34_005,inst_dob_i34_004,inst_dob_i34_003,inst_dob_i34_002,inst_dob_i34_001,inst_dob_i34_000}));
  // address_offset=18432;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_018432_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_Naddr_o_al_n54,addra[11:10]}),
    .csb({and_Naddrb$12$_Naddr_o_al_n57,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i36_008,inst_dob_i36_007,inst_dob_i36_006,inst_dob_i36_005,inst_dob_i36_004,inst_dob_i36_003,inst_dob_i36_002,inst_dob_i36_001,inst_dob_i36_000}));
  // address_offset=19456;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_019456_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_Naddr_o_al_n54,addra[11:10]}),
    .csb({and_Naddrb$12$_Naddr_o_al_n57,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i38_008,inst_dob_i38_007,inst_dob_i38_006,inst_dob_i38_005,inst_dob_i38_004,inst_dob_i38_003,inst_dob_i38_002,inst_dob_i38_001,inst_dob_i38_000}));
  // address_offset=20480;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_020480_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_Naddra_o_al_n70,addra[11:10]}),
    .csb({and_addrb$12$_Naddrb_o_al_n73,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i40_008,inst_dob_i40_007,inst_dob_i40_006,inst_dob_i40_005,inst_dob_i40_004,inst_dob_i40_003,inst_dob_i40_002,inst_dob_i40_001,inst_dob_i40_000}));
  // address_offset=21504;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_021504_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_Naddra_o_al_n70,addra[11:10]}),
    .csb({and_addrb$12$_Naddrb_o_al_n73,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i42_008,inst_dob_i42_007,inst_dob_i42_006,inst_dob_i42_005,inst_dob_i42_004,inst_dob_i42_003,inst_dob_i42_002,inst_dob_i42_001,inst_dob_i42_000}));
  // address_offset=22528;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_022528_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_Naddra_o_al_n70,addra[11:10]}),
    .csb({and_addrb$12$_Naddrb_o_al_n73,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i44_008,inst_dob_i44_007,inst_dob_i44_006,inst_dob_i44_005,inst_dob_i44_004,inst_dob_i44_003,inst_dob_i44_002,inst_dob_i44_001,inst_dob_i44_000}));
  // address_offset=23552;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_023552_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_Naddra_o_al_n70,addra[11:10]}),
    .csb({and_addrb$12$_Naddrb_o_al_n73,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i46_008,inst_dob_i46_007,inst_dob_i46_006,inst_dob_i46_005,inst_dob_i46_004,inst_dob_i46_003,inst_dob_i46_002,inst_dob_i46_001,inst_dob_i46_000}));
  // address_offset=24576;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_addra_o_al_n86,addra[11:10]}),
    .csb({and_Naddrb$12$_addrb_o_al_n89,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i48_008,inst_dob_i48_007,inst_dob_i48_006,inst_dob_i48_005,inst_dob_i48_004,inst_dob_i48_003,inst_dob_i48_002,inst_dob_i48_001,inst_dob_i48_000}));
  // address_offset=24576;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_009 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1395,open_n1396,open_n1397,open_n1398,open_n1399,open_n1400,open_n1401,dia[9],open_n1402}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1425,open_n1426,open_n1427,open_n1428,open_n1429,open_n1430,open_n1431,open_n1432,inst_dob_i48_009}));
  // address_offset=24576;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_010 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1433,open_n1434,open_n1435,open_n1436,open_n1437,open_n1438,open_n1439,dia[10],open_n1440}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1463,open_n1464,open_n1465,open_n1466,open_n1467,open_n1468,open_n1469,open_n1470,inst_dob_i48_010}));
  // address_offset=24576;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_011 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1471,open_n1472,open_n1473,open_n1474,open_n1475,open_n1476,open_n1477,dia[11],open_n1478}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1501,open_n1502,open_n1503,open_n1504,open_n1505,open_n1506,open_n1507,open_n1508,inst_dob_i48_011}));
  // address_offset=24576;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_012 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1509,open_n1510,open_n1511,open_n1512,open_n1513,open_n1514,open_n1515,dia[12],open_n1516}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1539,open_n1540,open_n1541,open_n1542,open_n1543,open_n1544,open_n1545,open_n1546,inst_dob_i48_012}));
  // address_offset=24576;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_013 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1547,open_n1548,open_n1549,open_n1550,open_n1551,open_n1552,open_n1553,dia[13],open_n1554}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1577,open_n1578,open_n1579,open_n1580,open_n1581,open_n1582,open_n1583,open_n1584,inst_dob_i48_013}));
  // address_offset=24576;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_014 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1585,open_n1586,open_n1587,open_n1588,open_n1589,open_n1590,open_n1591,dia[14],open_n1592}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1615,open_n1616,open_n1617,open_n1618,open_n1619,open_n1620,open_n1621,open_n1622,inst_dob_i48_014}));
  // address_offset=24576;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_015 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1623,open_n1624,open_n1625,open_n1626,open_n1627,open_n1628,open_n1629,dia[15],open_n1630}),
    .rsta(rsta),
    .rstb(rstb),
    .dob({open_n1653,open_n1654,open_n1655,open_n1656,open_n1657,open_n1658,open_n1659,open_n1660,inst_dob_i48_015}));
  // address_offset=25600;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_025600_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_addra_o_al_n86,addra[11:10]}),
    .csb({and_Naddrb$12$_addrb_o_al_n89,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i50_008,inst_dob_i50_007,inst_dob_i50_006,inst_dob_i50_005,inst_dob_i50_004,inst_dob_i50_003,inst_dob_i50_002,inst_dob_i50_001,inst_dob_i50_000}));
  // address_offset=26624;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_026624_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_addra_o_al_n86,addra[11:10]}),
    .csb({and_Naddrb$12$_addrb_o_al_n89,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i52_008,inst_dob_i52_007,inst_dob_i52_006,inst_dob_i52_005,inst_dob_i52_004,inst_dob_i52_003,inst_dob_i52_002,inst_dob_i52_001,inst_dob_i52_000}));
  // address_offset=27648;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_027648_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$12$_addra_o_al_n86,addra[11:10]}),
    .csb({and_Naddrb$12$_addrb_o_al_n89,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i54_008,inst_dob_i54_007,inst_dob_i54_006,inst_dob_i54_005,inst_dob_i54_004,inst_dob_i54_003,inst_dob_i54_002,inst_dob_i54_001,inst_dob_i54_000}));
  // address_offset=28672;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_028672_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_addra$_o_al_n102,addra[11:10]}),
    .csb({and_addrb$12$_addrb$_o_al_n105,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i56_008,inst_dob_i56_007,inst_dob_i56_006,inst_dob_i56_005,inst_dob_i56_004,inst_dob_i56_003,inst_dob_i56_002,inst_dob_i56_001,inst_dob_i56_000}));
  // address_offset=29696;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_029696_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_addra$_o_al_n102,addra[11:10]}),
    .csb({and_addrb$12$_addrb$_o_al_n105,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i58_008,inst_dob_i58_007,inst_dob_i58_006,inst_dob_i58_005,inst_dob_i58_004,inst_dob_i58_003,inst_dob_i58_002,inst_dob_i58_001,inst_dob_i58_000}));
  // address_offset=30720;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_030720_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_addra$_o_al_n102,addra[11:10]}),
    .csb({and_addrb$12$_addrb$_o_al_n105,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i60_008,inst_dob_i60_007,inst_dob_i60_006,inst_dob_i60_005,inst_dob_i60_004,inst_dob_i60_003,inst_dob_i60_002,inst_dob_i60_001,inst_dob_i60_000}));
  // address_offset=31744;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;address_step=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_031744_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({and_addra$12$_addra$_o_al_n102,addra[11:10]}),
    .csb({and_addrb$12$_addrb$_o_al_n105,addrb[11:10]}),
    .dia(dia[8:0]),
    .rsta(rsta),
    .rstb(rstb),
    .dob({inst_dob_i62_008,inst_dob_i62_007,inst_dob_i62_006,inst_dob_i62_005,inst_dob_i62_004,inst_dob_i62_003,inst_dob_i62_002,inst_dob_i62_001,inst_dob_i62_000}));
  // address_offset=32768;data_offset=0;depth=32;width=16;num_section=1;width_per_section=16;section_size=16;working_depth=512;working_width=18;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("18"),
    .DATA_WIDTH_B("18"),
    .MODE("PDPW8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_032768_000 (
    .addra({addra[8:0],4'b1111}),
    .addrb({addrb[8:0],4'b1111}),
    .clka(clka),
    .clkb(clkb),
    .csa({and_Naddra$11$_Naddr_o_and_cea,addra[10:9]}),
    .csb({and_Naddrb$11$_Naddr_o_and_ceb,addrb[10:9]}),
    .dia(dia[8:0]),
    .dib({open_n1817,open_n1818,dia[15:9]}),
    .rsta(rsta),
    .rstb(rstb),
    .doa({inst_dob_i64_008,inst_dob_i64_007,inst_dob_i64_006,inst_dob_i64_005,inst_dob_i64_004,inst_dob_i64_003,inst_dob_i64_002,inst_dob_i64_001,inst_dob_i64_000}),
    .dob({open_n1823,open_n1824,inst_dob_i64_015,inst_dob_i64_014,inst_dob_i64_013,inst_dob_i64_012,inst_dob_i64_011,inst_dob_i64_010,inst_dob_i64_009}));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_0  (
    .i0(inst_dob_i0_000),
    .i1(inst_dob_i0_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_1  (
    .i0(inst_dob_i2_000),
    .i1(inst_dob_i2_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_10  (
    .i0(inst_dob_i20_000),
    .i1(inst_dob_i20_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_10 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_11  (
    .i0(inst_dob_i22_000),
    .i1(inst_dob_i22_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_11 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_12  (
    .i0(inst_dob_i24_000),
    .i1(inst_dob_i24_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_12 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_13  (
    .i0(inst_dob_i26_000),
    .i1(inst_dob_i26_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_13 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_14  (
    .i0(inst_dob_i28_000),
    .i1(inst_dob_i28_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_14 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_15  (
    .i0(inst_dob_i30_000),
    .i1(inst_dob_i30_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_15 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_16  (
    .i0(inst_dob_i32_000),
    .i1(inst_dob_i32_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_16 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_17  (
    .i0(inst_dob_i34_000),
    .i1(inst_dob_i34_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_17 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_18  (
    .i0(inst_dob_i36_000),
    .i1(inst_dob_i36_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_18 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_19  (
    .i0(inst_dob_i38_000),
    .i1(inst_dob_i38_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_19 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_2  (
    .i0(inst_dob_i4_000),
    .i1(inst_dob_i4_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_20  (
    .i0(inst_dob_i40_000),
    .i1(inst_dob_i40_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_20 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_21  (
    .i0(inst_dob_i42_000),
    .i1(inst_dob_i42_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_21 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_22  (
    .i0(inst_dob_i44_000),
    .i1(inst_dob_i44_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_22 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_23  (
    .i0(inst_dob_i46_000),
    .i1(inst_dob_i46_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_23 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_24  (
    .i0(inst_dob_i48_000),
    .i1(inst_dob_i48_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_24 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_25  (
    .i0(inst_dob_i50_000),
    .i1(inst_dob_i50_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_25 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_26  (
    .i0(inst_dob_i52_000),
    .i1(inst_dob_i52_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_26 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_27  (
    .i0(inst_dob_i54_000),
    .i1(inst_dob_i54_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_27 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_28  (
    .i0(inst_dob_i56_000),
    .i1(inst_dob_i56_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_28 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_29  (
    .i0(inst_dob_i58_000),
    .i1(inst_dob_i58_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_29 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_3  (
    .i0(inst_dob_i6_000),
    .i1(inst_dob_i6_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_30  (
    .i0(inst_dob_i60_000),
    .i1(inst_dob_i60_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_30 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_31  (
    .i0(inst_dob_i62_000),
    .i1(inst_dob_i62_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_31 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_32  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_32 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_33  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_33 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_34  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_34 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_35  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_35 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_36  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_36 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_37  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_37 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_38  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_38 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_39  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_39 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_4  (
    .i0(inst_dob_i8_000),
    .i1(inst_dob_i8_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_4 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_40  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_40 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_41  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_41 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_42  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_42 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_43  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_43 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_44  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_44 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_45  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_45 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_46  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_46 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_47  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_47 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_48  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_48 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_49  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_49 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_5  (
    .i0(inst_dob_i10_000),
    .i1(inst_dob_i10_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_5 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_50  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_50 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_51  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_51 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_52  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_52 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_53  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_53 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_54  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_54 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_55  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_55 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_56  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_56 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_57  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_57 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_58  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_58 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_59  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_59 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_6  (
    .i0(inst_dob_i12_000),
    .i1(inst_dob_i12_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_6 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_60  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_60 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_61  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_61 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_62  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_62 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_63  (
    .i0(inst_dob_i64_000),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_63 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_7  (
    .i0(inst_dob_i14_000),
    .i1(inst_dob_i14_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_7 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_8  (
    .i0(inst_dob_i16_000),
    .i1(inst_dob_i16_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_8 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_9  (
    .i0(inst_dob_i18_000),
    .i1(inst_dob_i18_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_9 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b0/B0_0 ),
    .i1(\inst_dob_mux_b0/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b0/B0_2 ),
    .i1(\inst_dob_mux_b0/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b0/B0_20 ),
    .i1(\inst_dob_mux_b0/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_10 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b0/B0_22 ),
    .i1(\inst_dob_mux_b0/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_11 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b0/B0_24 ),
    .i1(\inst_dob_mux_b0/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_12 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b0/B0_26 ),
    .i1(\inst_dob_mux_b0/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_13 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b0/B0_28 ),
    .i1(\inst_dob_mux_b0/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_14 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b0/B0_30 ),
    .i1(\inst_dob_mux_b0/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_15 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b0/B0_32 ),
    .i1(\inst_dob_mux_b0/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_16 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b0/B0_34 ),
    .i1(\inst_dob_mux_b0/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_17 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b0/B0_36 ),
    .i1(\inst_dob_mux_b0/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_18 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b0/B0_38 ),
    .i1(\inst_dob_mux_b0/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_19 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b0/B0_4 ),
    .i1(\inst_dob_mux_b0/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b0/B0_40 ),
    .i1(\inst_dob_mux_b0/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_20 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b0/B0_42 ),
    .i1(\inst_dob_mux_b0/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_21 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b0/B0_44 ),
    .i1(\inst_dob_mux_b0/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_22 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b0/B0_46 ),
    .i1(\inst_dob_mux_b0/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_23 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b0/B0_48 ),
    .i1(\inst_dob_mux_b0/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_24 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b0/B0_50 ),
    .i1(\inst_dob_mux_b0/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_25 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b0/B0_52 ),
    .i1(\inst_dob_mux_b0/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_26 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b0/B0_54 ),
    .i1(\inst_dob_mux_b0/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_27 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b0/B0_56 ),
    .i1(\inst_dob_mux_b0/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_28 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b0/B0_58 ),
    .i1(\inst_dob_mux_b0/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_29 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b0/B0_6 ),
    .i1(\inst_dob_mux_b0/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b0/B0_60 ),
    .i1(\inst_dob_mux_b0/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_30 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b0/B0_62 ),
    .i1(\inst_dob_mux_b0/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_31 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b0/B0_8 ),
    .i1(\inst_dob_mux_b0/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_4 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b0/B0_10 ),
    .i1(\inst_dob_mux_b0/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_5 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b0/B0_12 ),
    .i1(\inst_dob_mux_b0/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_6 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b0/B0_14 ),
    .i1(\inst_dob_mux_b0/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_7 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b0/B0_16 ),
    .i1(\inst_dob_mux_b0/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_8 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b0/B0_18 ),
    .i1(\inst_dob_mux_b0/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_9 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b0/B1_0 ),
    .i1(\inst_dob_mux_b0/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b0/B1_2 ),
    .i1(\inst_dob_mux_b0/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b0/B1_20 ),
    .i1(\inst_dob_mux_b0/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_10 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b0/B1_22 ),
    .i1(\inst_dob_mux_b0/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_11 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b0/B1_24 ),
    .i1(\inst_dob_mux_b0/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_12 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b0/B1_26 ),
    .i1(\inst_dob_mux_b0/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_13 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b0/B1_28 ),
    .i1(\inst_dob_mux_b0/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_14 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b0/B1_30 ),
    .i1(\inst_dob_mux_b0/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_15 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b0/B1_4 ),
    .i1(\inst_dob_mux_b0/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b0/B1_6 ),
    .i1(\inst_dob_mux_b0/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b0/B1_8 ),
    .i1(\inst_dob_mux_b0/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_4 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b0/B1_10 ),
    .i1(\inst_dob_mux_b0/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_5 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b0/B1_12 ),
    .i1(\inst_dob_mux_b0/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_6 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b0/B1_14 ),
    .i1(\inst_dob_mux_b0/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_7 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b0/B1_16 ),
    .i1(\inst_dob_mux_b0/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_8 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b0/B1_18 ),
    .i1(\inst_dob_mux_b0/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_9 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b0/B2_0 ),
    .i1(\inst_dob_mux_b0/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b0/B3_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b0/B2_2 ),
    .i1(\inst_dob_mux_b0/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b0/B3_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b0/B2_4 ),
    .i1(\inst_dob_mux_b0/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b0/B3_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b0/B2_6 ),
    .i1(\inst_dob_mux_b0/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b0/B3_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b0/B2_8 ),
    .i1(\inst_dob_mux_b0/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b0/B3_4 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b0/B2_10 ),
    .i1(\inst_dob_mux_b0/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b0/B3_5 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b0/B2_12 ),
    .i1(\inst_dob_mux_b0/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b0/B3_6 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b0/B2_14 ),
    .i1(\inst_dob_mux_b0/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b0/B3_7 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b0/B3_0 ),
    .i1(\inst_dob_mux_b0/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b0/B4_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b0/B3_2 ),
    .i1(\inst_dob_mux_b0/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b0/B4_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b0/B3_4 ),
    .i1(\inst_dob_mux_b0/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b0/B4_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b0/B3_6 ),
    .i1(\inst_dob_mux_b0/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b0/B4_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b0/B4_0 ),
    .i1(\inst_dob_mux_b0/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b0/B5_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b0/B4_2 ),
    .i1(\inst_dob_mux_b0/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b0/B5_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b0/B5_0 ),
    .i1(\inst_dob_mux_b0/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[0]));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_0  (
    .i0(inst_dob_i0_001),
    .i1(inst_dob_i0_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_1  (
    .i0(inst_dob_i2_001),
    .i1(inst_dob_i2_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_10  (
    .i0(inst_dob_i20_001),
    .i1(inst_dob_i20_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_10 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_11  (
    .i0(inst_dob_i22_001),
    .i1(inst_dob_i22_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_11 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_12  (
    .i0(inst_dob_i24_001),
    .i1(inst_dob_i24_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_12 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_13  (
    .i0(inst_dob_i26_001),
    .i1(inst_dob_i26_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_13 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_14  (
    .i0(inst_dob_i28_001),
    .i1(inst_dob_i28_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_14 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_15  (
    .i0(inst_dob_i30_001),
    .i1(inst_dob_i30_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_15 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_16  (
    .i0(inst_dob_i32_001),
    .i1(inst_dob_i32_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_16 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_17  (
    .i0(inst_dob_i34_001),
    .i1(inst_dob_i34_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_17 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_18  (
    .i0(inst_dob_i36_001),
    .i1(inst_dob_i36_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_18 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_19  (
    .i0(inst_dob_i38_001),
    .i1(inst_dob_i38_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_19 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_2  (
    .i0(inst_dob_i4_001),
    .i1(inst_dob_i4_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_20  (
    .i0(inst_dob_i40_001),
    .i1(inst_dob_i40_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_20 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_21  (
    .i0(inst_dob_i42_001),
    .i1(inst_dob_i42_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_21 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_22  (
    .i0(inst_dob_i44_001),
    .i1(inst_dob_i44_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_22 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_23  (
    .i0(inst_dob_i46_001),
    .i1(inst_dob_i46_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_23 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_24  (
    .i0(inst_dob_i48_001),
    .i1(inst_dob_i48_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_24 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_25  (
    .i0(inst_dob_i50_001),
    .i1(inst_dob_i50_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_25 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_26  (
    .i0(inst_dob_i52_001),
    .i1(inst_dob_i52_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_26 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_27  (
    .i0(inst_dob_i54_001),
    .i1(inst_dob_i54_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_27 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_28  (
    .i0(inst_dob_i56_001),
    .i1(inst_dob_i56_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_28 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_29  (
    .i0(inst_dob_i58_001),
    .i1(inst_dob_i58_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_29 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_3  (
    .i0(inst_dob_i6_001),
    .i1(inst_dob_i6_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_30  (
    .i0(inst_dob_i60_001),
    .i1(inst_dob_i60_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_30 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_31  (
    .i0(inst_dob_i62_001),
    .i1(inst_dob_i62_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_31 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_32  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_32 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_33  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_33 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_34  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_34 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_35  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_35 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_36  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_36 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_37  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_37 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_38  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_38 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_39  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_39 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_4  (
    .i0(inst_dob_i8_001),
    .i1(inst_dob_i8_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_4 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_40  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_40 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_41  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_41 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_42  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_42 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_43  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_43 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_44  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_44 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_45  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_45 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_46  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_46 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_47  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_47 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_48  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_48 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_49  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_49 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_5  (
    .i0(inst_dob_i10_001),
    .i1(inst_dob_i10_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_5 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_50  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_50 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_51  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_51 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_52  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_52 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_53  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_53 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_54  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_54 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_55  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_55 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_56  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_56 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_57  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_57 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_58  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_58 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_59  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_59 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_6  (
    .i0(inst_dob_i12_001),
    .i1(inst_dob_i12_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_6 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_60  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_60 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_61  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_61 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_62  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_62 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_63  (
    .i0(inst_dob_i64_001),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_63 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_7  (
    .i0(inst_dob_i14_001),
    .i1(inst_dob_i14_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_7 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_8  (
    .i0(inst_dob_i16_001),
    .i1(inst_dob_i16_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_8 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_9  (
    .i0(inst_dob_i18_001),
    .i1(inst_dob_i18_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_9 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b1/B0_0 ),
    .i1(\inst_dob_mux_b1/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b1/B0_2 ),
    .i1(\inst_dob_mux_b1/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b1/B0_20 ),
    .i1(\inst_dob_mux_b1/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_10 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b1/B0_22 ),
    .i1(\inst_dob_mux_b1/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_11 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b1/B0_24 ),
    .i1(\inst_dob_mux_b1/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_12 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b1/B0_26 ),
    .i1(\inst_dob_mux_b1/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_13 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b1/B0_28 ),
    .i1(\inst_dob_mux_b1/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_14 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b1/B0_30 ),
    .i1(\inst_dob_mux_b1/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_15 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b1/B0_32 ),
    .i1(\inst_dob_mux_b1/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_16 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b1/B0_34 ),
    .i1(\inst_dob_mux_b1/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_17 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b1/B0_36 ),
    .i1(\inst_dob_mux_b1/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_18 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b1/B0_38 ),
    .i1(\inst_dob_mux_b1/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_19 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b1/B0_4 ),
    .i1(\inst_dob_mux_b1/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b1/B0_40 ),
    .i1(\inst_dob_mux_b1/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_20 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b1/B0_42 ),
    .i1(\inst_dob_mux_b1/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_21 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b1/B0_44 ),
    .i1(\inst_dob_mux_b1/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_22 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b1/B0_46 ),
    .i1(\inst_dob_mux_b1/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_23 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b1/B0_48 ),
    .i1(\inst_dob_mux_b1/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_24 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b1/B0_50 ),
    .i1(\inst_dob_mux_b1/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_25 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b1/B0_52 ),
    .i1(\inst_dob_mux_b1/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_26 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b1/B0_54 ),
    .i1(\inst_dob_mux_b1/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_27 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b1/B0_56 ),
    .i1(\inst_dob_mux_b1/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_28 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b1/B0_58 ),
    .i1(\inst_dob_mux_b1/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_29 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b1/B0_6 ),
    .i1(\inst_dob_mux_b1/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b1/B0_60 ),
    .i1(\inst_dob_mux_b1/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_30 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b1/B0_62 ),
    .i1(\inst_dob_mux_b1/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_31 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b1/B0_8 ),
    .i1(\inst_dob_mux_b1/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_4 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b1/B0_10 ),
    .i1(\inst_dob_mux_b1/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_5 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b1/B0_12 ),
    .i1(\inst_dob_mux_b1/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_6 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b1/B0_14 ),
    .i1(\inst_dob_mux_b1/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_7 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b1/B0_16 ),
    .i1(\inst_dob_mux_b1/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_8 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b1/B0_18 ),
    .i1(\inst_dob_mux_b1/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_9 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b1/B1_0 ),
    .i1(\inst_dob_mux_b1/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b1/B1_2 ),
    .i1(\inst_dob_mux_b1/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b1/B1_20 ),
    .i1(\inst_dob_mux_b1/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_10 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b1/B1_22 ),
    .i1(\inst_dob_mux_b1/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_11 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b1/B1_24 ),
    .i1(\inst_dob_mux_b1/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_12 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b1/B1_26 ),
    .i1(\inst_dob_mux_b1/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_13 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b1/B1_28 ),
    .i1(\inst_dob_mux_b1/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_14 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b1/B1_30 ),
    .i1(\inst_dob_mux_b1/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_15 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b1/B1_4 ),
    .i1(\inst_dob_mux_b1/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b1/B1_6 ),
    .i1(\inst_dob_mux_b1/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b1/B1_8 ),
    .i1(\inst_dob_mux_b1/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_4 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b1/B1_10 ),
    .i1(\inst_dob_mux_b1/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_5 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b1/B1_12 ),
    .i1(\inst_dob_mux_b1/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_6 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b1/B1_14 ),
    .i1(\inst_dob_mux_b1/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_7 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b1/B1_16 ),
    .i1(\inst_dob_mux_b1/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_8 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b1/B1_18 ),
    .i1(\inst_dob_mux_b1/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_9 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b1/B2_0 ),
    .i1(\inst_dob_mux_b1/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b1/B3_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b1/B2_2 ),
    .i1(\inst_dob_mux_b1/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b1/B3_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b1/B2_4 ),
    .i1(\inst_dob_mux_b1/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b1/B3_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b1/B2_6 ),
    .i1(\inst_dob_mux_b1/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b1/B3_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b1/B2_8 ),
    .i1(\inst_dob_mux_b1/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b1/B3_4 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b1/B2_10 ),
    .i1(\inst_dob_mux_b1/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b1/B3_5 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b1/B2_12 ),
    .i1(\inst_dob_mux_b1/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b1/B3_6 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b1/B2_14 ),
    .i1(\inst_dob_mux_b1/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b1/B3_7 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b1/B3_0 ),
    .i1(\inst_dob_mux_b1/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b1/B4_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b1/B3_2 ),
    .i1(\inst_dob_mux_b1/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b1/B4_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b1/B3_4 ),
    .i1(\inst_dob_mux_b1/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b1/B4_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b1/B3_6 ),
    .i1(\inst_dob_mux_b1/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b1/B4_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b1/B4_0 ),
    .i1(\inst_dob_mux_b1/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b1/B5_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b1/B4_2 ),
    .i1(\inst_dob_mux_b1/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b1/B5_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b1/B5_0 ),
    .i1(\inst_dob_mux_b1/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[1]));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_0  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_1  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_10  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_10 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_11  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_11 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_12  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_12 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_13  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_13 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_14  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_14 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_15  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_15 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_16  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_16 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_17  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_17 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_18  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_18 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_19  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_19 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_2  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_2 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_20  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_20 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_21  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_21 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_22  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_22 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_23  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i32_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_23 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_24  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_24 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_25  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_25 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_26  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_26 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_27  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_27 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_28  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_28 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_29  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_29 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_3  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_3 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_30  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_30 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_31  (
    .i0(inst_dob_i48_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_31 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_32  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_32 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_33  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_33 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_34  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_34 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_35  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_35 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_36  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_36 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_37  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_37 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_38  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_38 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_39  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_39 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_4  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_4 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_40  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_40 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_41  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_41 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_42  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_42 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_43  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_43 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_44  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_44 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_45  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_45 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_46  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_46 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_47  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_47 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_48  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_48 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_49  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_49 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_5  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_5 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_50  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_50 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_51  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_51 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_52  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_52 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_53  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_53 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_54  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_54 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_55  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_55 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_56  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_56 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_57  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_57 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_58  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_58 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_59  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_59 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_6  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_6 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_60  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_60 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_61  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_61 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_62  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_62 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_63  (
    .i0(inst_dob_i64_010),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_63 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_7  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i0_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_7 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_8  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_8 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_9  (
    .i0(inst_dob_i16_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_9 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b10/B0_0 ),
    .i1(\inst_dob_mux_b10/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b10/B0_2 ),
    .i1(\inst_dob_mux_b10/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b10/B0_20 ),
    .i1(\inst_dob_mux_b10/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_10 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b10/B0_22 ),
    .i1(\inst_dob_mux_b10/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_11 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b10/B0_24 ),
    .i1(\inst_dob_mux_b10/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_12 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b10/B0_26 ),
    .i1(\inst_dob_mux_b10/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_13 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b10/B0_28 ),
    .i1(\inst_dob_mux_b10/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_14 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b10/B0_30 ),
    .i1(\inst_dob_mux_b10/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_15 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b10/B0_32 ),
    .i1(\inst_dob_mux_b10/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_16 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b10/B0_34 ),
    .i1(\inst_dob_mux_b10/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_17 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b10/B0_36 ),
    .i1(\inst_dob_mux_b10/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_18 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b10/B0_38 ),
    .i1(\inst_dob_mux_b10/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_19 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b10/B0_4 ),
    .i1(\inst_dob_mux_b10/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_2 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b10/B0_40 ),
    .i1(\inst_dob_mux_b10/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_20 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b10/B0_42 ),
    .i1(\inst_dob_mux_b10/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_21 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b10/B0_44 ),
    .i1(\inst_dob_mux_b10/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_22 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b10/B0_46 ),
    .i1(\inst_dob_mux_b10/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_23 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b10/B0_48 ),
    .i1(\inst_dob_mux_b10/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_24 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b10/B0_50 ),
    .i1(\inst_dob_mux_b10/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_25 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b10/B0_52 ),
    .i1(\inst_dob_mux_b10/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_26 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b10/B0_54 ),
    .i1(\inst_dob_mux_b10/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_27 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b10/B0_56 ),
    .i1(\inst_dob_mux_b10/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_28 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b10/B0_58 ),
    .i1(\inst_dob_mux_b10/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_29 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b10/B0_6 ),
    .i1(\inst_dob_mux_b10/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_3 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b10/B0_60 ),
    .i1(\inst_dob_mux_b10/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_30 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b10/B0_62 ),
    .i1(\inst_dob_mux_b10/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_31 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b10/B0_8 ),
    .i1(\inst_dob_mux_b10/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_4 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b10/B0_10 ),
    .i1(\inst_dob_mux_b10/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_5 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b10/B0_12 ),
    .i1(\inst_dob_mux_b10/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_6 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b10/B0_14 ),
    .i1(\inst_dob_mux_b10/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_7 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b10/B0_16 ),
    .i1(\inst_dob_mux_b10/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_8 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b10/B0_18 ),
    .i1(\inst_dob_mux_b10/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_9 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b10/B1_0 ),
    .i1(\inst_dob_mux_b10/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b10/B1_2 ),
    .i1(\inst_dob_mux_b10/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b10/B1_20 ),
    .i1(\inst_dob_mux_b10/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_10 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b10/B1_22 ),
    .i1(\inst_dob_mux_b10/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_11 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b10/B1_24 ),
    .i1(\inst_dob_mux_b10/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_12 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b10/B1_26 ),
    .i1(\inst_dob_mux_b10/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_13 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b10/B1_28 ),
    .i1(\inst_dob_mux_b10/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_14 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b10/B1_30 ),
    .i1(\inst_dob_mux_b10/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_15 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b10/B1_4 ),
    .i1(\inst_dob_mux_b10/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_2 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b10/B1_6 ),
    .i1(\inst_dob_mux_b10/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_3 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b10/B1_8 ),
    .i1(\inst_dob_mux_b10/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_4 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b10/B1_10 ),
    .i1(\inst_dob_mux_b10/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_5 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b10/B1_12 ),
    .i1(\inst_dob_mux_b10/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_6 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b10/B1_14 ),
    .i1(\inst_dob_mux_b10/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_7 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b10/B1_16 ),
    .i1(\inst_dob_mux_b10/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_8 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b10/B1_18 ),
    .i1(\inst_dob_mux_b10/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b10/B2_9 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b10/B2_0 ),
    .i1(\inst_dob_mux_b10/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b10/B3_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b10/B2_2 ),
    .i1(\inst_dob_mux_b10/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b10/B3_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b10/B2_4 ),
    .i1(\inst_dob_mux_b10/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b10/B3_2 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b10/B2_6 ),
    .i1(\inst_dob_mux_b10/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b10/B3_3 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b10/B2_8 ),
    .i1(\inst_dob_mux_b10/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b10/B3_4 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b10/B2_10 ),
    .i1(\inst_dob_mux_b10/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b10/B3_5 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b10/B2_12 ),
    .i1(\inst_dob_mux_b10/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b10/B3_6 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b10/B2_14 ),
    .i1(\inst_dob_mux_b10/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b10/B3_7 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b10/B3_0 ),
    .i1(\inst_dob_mux_b10/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b10/B4_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b10/B3_2 ),
    .i1(\inst_dob_mux_b10/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b10/B4_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b10/B3_4 ),
    .i1(\inst_dob_mux_b10/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b10/B4_2 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b10/B3_6 ),
    .i1(\inst_dob_mux_b10/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b10/B4_3 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b10/B4_0 ),
    .i1(\inst_dob_mux_b10/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b10/B5_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b10/B4_2 ),
    .i1(\inst_dob_mux_b10/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b10/B5_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b10/B5_0 ),
    .i1(\inst_dob_mux_b10/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[10]));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_0  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_1  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_10  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_10 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_11  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_11 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_12  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_12 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_13  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_13 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_14  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_14 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_15  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_15 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_16  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_16 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_17  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_17 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_18  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_18 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_19  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_19 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_2  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_2 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_20  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_20 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_21  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_21 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_22  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_22 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_23  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i32_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_23 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_24  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_24 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_25  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_25 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_26  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_26 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_27  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_27 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_28  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_28 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_29  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_29 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_3  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_3 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_30  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_30 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_31  (
    .i0(inst_dob_i48_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_31 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_32  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_32 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_33  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_33 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_34  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_34 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_35  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_35 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_36  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_36 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_37  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_37 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_38  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_38 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_39  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_39 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_4  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_4 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_40  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_40 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_41  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_41 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_42  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_42 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_43  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_43 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_44  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_44 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_45  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_45 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_46  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_46 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_47  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_47 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_48  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_48 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_49  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_49 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_5  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_5 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_50  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_50 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_51  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_51 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_52  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_52 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_53  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_53 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_54  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_54 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_55  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_55 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_56  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_56 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_57  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_57 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_58  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_58 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_59  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_59 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_6  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_6 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_60  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_60 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_61  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_61 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_62  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_62 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_63  (
    .i0(inst_dob_i64_011),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_63 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_7  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i0_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_7 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_8  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_8 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_9  (
    .i0(inst_dob_i16_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_9 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b11/B0_0 ),
    .i1(\inst_dob_mux_b11/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b11/B0_2 ),
    .i1(\inst_dob_mux_b11/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b11/B0_20 ),
    .i1(\inst_dob_mux_b11/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_10 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b11/B0_22 ),
    .i1(\inst_dob_mux_b11/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_11 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b11/B0_24 ),
    .i1(\inst_dob_mux_b11/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_12 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b11/B0_26 ),
    .i1(\inst_dob_mux_b11/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_13 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b11/B0_28 ),
    .i1(\inst_dob_mux_b11/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_14 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b11/B0_30 ),
    .i1(\inst_dob_mux_b11/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_15 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b11/B0_32 ),
    .i1(\inst_dob_mux_b11/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_16 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b11/B0_34 ),
    .i1(\inst_dob_mux_b11/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_17 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b11/B0_36 ),
    .i1(\inst_dob_mux_b11/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_18 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b11/B0_38 ),
    .i1(\inst_dob_mux_b11/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_19 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b11/B0_4 ),
    .i1(\inst_dob_mux_b11/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_2 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b11/B0_40 ),
    .i1(\inst_dob_mux_b11/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_20 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b11/B0_42 ),
    .i1(\inst_dob_mux_b11/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_21 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b11/B0_44 ),
    .i1(\inst_dob_mux_b11/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_22 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b11/B0_46 ),
    .i1(\inst_dob_mux_b11/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_23 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b11/B0_48 ),
    .i1(\inst_dob_mux_b11/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_24 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b11/B0_50 ),
    .i1(\inst_dob_mux_b11/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_25 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b11/B0_52 ),
    .i1(\inst_dob_mux_b11/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_26 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b11/B0_54 ),
    .i1(\inst_dob_mux_b11/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_27 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b11/B0_56 ),
    .i1(\inst_dob_mux_b11/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_28 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b11/B0_58 ),
    .i1(\inst_dob_mux_b11/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_29 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b11/B0_6 ),
    .i1(\inst_dob_mux_b11/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_3 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b11/B0_60 ),
    .i1(\inst_dob_mux_b11/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_30 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b11/B0_62 ),
    .i1(\inst_dob_mux_b11/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_31 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b11/B0_8 ),
    .i1(\inst_dob_mux_b11/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_4 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b11/B0_10 ),
    .i1(\inst_dob_mux_b11/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_5 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b11/B0_12 ),
    .i1(\inst_dob_mux_b11/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_6 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b11/B0_14 ),
    .i1(\inst_dob_mux_b11/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_7 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b11/B0_16 ),
    .i1(\inst_dob_mux_b11/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_8 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b11/B0_18 ),
    .i1(\inst_dob_mux_b11/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_9 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b11/B1_0 ),
    .i1(\inst_dob_mux_b11/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b11/B1_2 ),
    .i1(\inst_dob_mux_b11/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b11/B1_20 ),
    .i1(\inst_dob_mux_b11/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_10 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b11/B1_22 ),
    .i1(\inst_dob_mux_b11/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_11 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b11/B1_24 ),
    .i1(\inst_dob_mux_b11/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_12 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b11/B1_26 ),
    .i1(\inst_dob_mux_b11/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_13 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b11/B1_28 ),
    .i1(\inst_dob_mux_b11/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_14 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b11/B1_30 ),
    .i1(\inst_dob_mux_b11/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_15 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b11/B1_4 ),
    .i1(\inst_dob_mux_b11/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_2 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b11/B1_6 ),
    .i1(\inst_dob_mux_b11/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_3 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b11/B1_8 ),
    .i1(\inst_dob_mux_b11/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_4 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b11/B1_10 ),
    .i1(\inst_dob_mux_b11/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_5 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b11/B1_12 ),
    .i1(\inst_dob_mux_b11/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_6 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b11/B1_14 ),
    .i1(\inst_dob_mux_b11/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_7 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b11/B1_16 ),
    .i1(\inst_dob_mux_b11/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_8 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b11/B1_18 ),
    .i1(\inst_dob_mux_b11/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b11/B2_9 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b11/B2_0 ),
    .i1(\inst_dob_mux_b11/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b11/B3_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b11/B2_2 ),
    .i1(\inst_dob_mux_b11/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b11/B3_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b11/B2_4 ),
    .i1(\inst_dob_mux_b11/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b11/B3_2 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b11/B2_6 ),
    .i1(\inst_dob_mux_b11/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b11/B3_3 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b11/B2_8 ),
    .i1(\inst_dob_mux_b11/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b11/B3_4 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b11/B2_10 ),
    .i1(\inst_dob_mux_b11/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b11/B3_5 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b11/B2_12 ),
    .i1(\inst_dob_mux_b11/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b11/B3_6 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b11/B2_14 ),
    .i1(\inst_dob_mux_b11/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b11/B3_7 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b11/B3_0 ),
    .i1(\inst_dob_mux_b11/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b11/B4_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b11/B3_2 ),
    .i1(\inst_dob_mux_b11/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b11/B4_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b11/B3_4 ),
    .i1(\inst_dob_mux_b11/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b11/B4_2 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b11/B3_6 ),
    .i1(\inst_dob_mux_b11/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b11/B4_3 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b11/B4_0 ),
    .i1(\inst_dob_mux_b11/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b11/B5_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b11/B4_2 ),
    .i1(\inst_dob_mux_b11/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b11/B5_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b11/B5_0 ),
    .i1(\inst_dob_mux_b11/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[11]));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_0  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_1  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_10  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_10 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_11  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_11 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_12  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_12 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_13  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_13 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_14  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_14 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_15  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_15 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_16  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_16 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_17  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_17 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_18  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_18 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_19  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_19 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_2  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_2 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_20  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_20 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_21  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_21 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_22  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_22 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_23  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i32_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_23 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_24  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_24 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_25  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_25 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_26  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_26 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_27  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_27 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_28  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_28 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_29  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_29 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_3  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_3 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_30  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_30 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_31  (
    .i0(inst_dob_i48_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_31 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_32  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_32 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_33  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_33 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_34  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_34 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_35  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_35 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_36  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_36 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_37  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_37 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_38  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_38 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_39  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_39 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_4  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_4 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_40  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_40 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_41  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_41 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_42  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_42 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_43  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_43 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_44  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_44 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_45  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_45 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_46  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_46 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_47  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_47 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_48  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_48 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_49  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_49 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_5  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_5 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_50  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_50 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_51  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_51 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_52  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_52 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_53  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_53 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_54  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_54 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_55  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_55 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_56  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_56 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_57  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_57 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_58  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_58 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_59  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_59 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_6  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_6 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_60  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_60 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_61  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_61 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_62  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_62 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_63  (
    .i0(inst_dob_i64_012),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_63 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_7  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i0_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_7 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_8  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_8 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_9  (
    .i0(inst_dob_i16_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_9 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b12/B0_0 ),
    .i1(\inst_dob_mux_b12/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b12/B0_2 ),
    .i1(\inst_dob_mux_b12/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b12/B0_20 ),
    .i1(\inst_dob_mux_b12/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_10 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b12/B0_22 ),
    .i1(\inst_dob_mux_b12/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_11 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b12/B0_24 ),
    .i1(\inst_dob_mux_b12/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_12 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b12/B0_26 ),
    .i1(\inst_dob_mux_b12/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_13 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b12/B0_28 ),
    .i1(\inst_dob_mux_b12/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_14 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b12/B0_30 ),
    .i1(\inst_dob_mux_b12/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_15 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b12/B0_32 ),
    .i1(\inst_dob_mux_b12/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_16 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b12/B0_34 ),
    .i1(\inst_dob_mux_b12/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_17 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b12/B0_36 ),
    .i1(\inst_dob_mux_b12/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_18 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b12/B0_38 ),
    .i1(\inst_dob_mux_b12/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_19 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b12/B0_4 ),
    .i1(\inst_dob_mux_b12/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_2 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b12/B0_40 ),
    .i1(\inst_dob_mux_b12/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_20 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b12/B0_42 ),
    .i1(\inst_dob_mux_b12/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_21 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b12/B0_44 ),
    .i1(\inst_dob_mux_b12/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_22 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b12/B0_46 ),
    .i1(\inst_dob_mux_b12/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_23 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b12/B0_48 ),
    .i1(\inst_dob_mux_b12/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_24 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b12/B0_50 ),
    .i1(\inst_dob_mux_b12/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_25 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b12/B0_52 ),
    .i1(\inst_dob_mux_b12/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_26 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b12/B0_54 ),
    .i1(\inst_dob_mux_b12/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_27 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b12/B0_56 ),
    .i1(\inst_dob_mux_b12/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_28 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b12/B0_58 ),
    .i1(\inst_dob_mux_b12/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_29 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b12/B0_6 ),
    .i1(\inst_dob_mux_b12/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_3 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b12/B0_60 ),
    .i1(\inst_dob_mux_b12/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_30 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b12/B0_62 ),
    .i1(\inst_dob_mux_b12/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_31 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b12/B0_8 ),
    .i1(\inst_dob_mux_b12/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_4 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b12/B0_10 ),
    .i1(\inst_dob_mux_b12/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_5 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b12/B0_12 ),
    .i1(\inst_dob_mux_b12/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_6 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b12/B0_14 ),
    .i1(\inst_dob_mux_b12/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_7 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b12/B0_16 ),
    .i1(\inst_dob_mux_b12/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_8 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b12/B0_18 ),
    .i1(\inst_dob_mux_b12/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_9 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b12/B1_0 ),
    .i1(\inst_dob_mux_b12/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b12/B1_2 ),
    .i1(\inst_dob_mux_b12/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b12/B1_20 ),
    .i1(\inst_dob_mux_b12/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_10 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b12/B1_22 ),
    .i1(\inst_dob_mux_b12/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_11 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b12/B1_24 ),
    .i1(\inst_dob_mux_b12/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_12 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b12/B1_26 ),
    .i1(\inst_dob_mux_b12/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_13 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b12/B1_28 ),
    .i1(\inst_dob_mux_b12/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_14 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b12/B1_30 ),
    .i1(\inst_dob_mux_b12/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_15 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b12/B1_4 ),
    .i1(\inst_dob_mux_b12/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_2 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b12/B1_6 ),
    .i1(\inst_dob_mux_b12/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_3 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b12/B1_8 ),
    .i1(\inst_dob_mux_b12/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_4 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b12/B1_10 ),
    .i1(\inst_dob_mux_b12/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_5 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b12/B1_12 ),
    .i1(\inst_dob_mux_b12/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_6 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b12/B1_14 ),
    .i1(\inst_dob_mux_b12/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_7 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b12/B1_16 ),
    .i1(\inst_dob_mux_b12/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_8 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b12/B1_18 ),
    .i1(\inst_dob_mux_b12/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b12/B2_9 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b12/B2_0 ),
    .i1(\inst_dob_mux_b12/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b12/B3_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b12/B2_2 ),
    .i1(\inst_dob_mux_b12/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b12/B3_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b12/B2_4 ),
    .i1(\inst_dob_mux_b12/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b12/B3_2 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b12/B2_6 ),
    .i1(\inst_dob_mux_b12/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b12/B3_3 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b12/B2_8 ),
    .i1(\inst_dob_mux_b12/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b12/B3_4 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b12/B2_10 ),
    .i1(\inst_dob_mux_b12/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b12/B3_5 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b12/B2_12 ),
    .i1(\inst_dob_mux_b12/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b12/B3_6 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b12/B2_14 ),
    .i1(\inst_dob_mux_b12/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b12/B3_7 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b12/B3_0 ),
    .i1(\inst_dob_mux_b12/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b12/B4_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b12/B3_2 ),
    .i1(\inst_dob_mux_b12/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b12/B4_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b12/B3_4 ),
    .i1(\inst_dob_mux_b12/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b12/B4_2 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b12/B3_6 ),
    .i1(\inst_dob_mux_b12/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b12/B4_3 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b12/B4_0 ),
    .i1(\inst_dob_mux_b12/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b12/B5_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b12/B4_2 ),
    .i1(\inst_dob_mux_b12/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b12/B5_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b12/B5_0 ),
    .i1(\inst_dob_mux_b12/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[12]));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_0  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_1  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_10  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_10 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_11  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_11 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_12  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_12 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_13  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_13 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_14  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_14 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_15  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_15 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_16  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_16 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_17  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_17 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_18  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_18 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_19  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_19 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_2  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_2 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_20  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_20 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_21  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_21 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_22  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_22 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_23  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i32_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_23 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_24  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_24 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_25  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_25 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_26  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_26 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_27  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_27 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_28  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_28 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_29  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_29 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_3  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_3 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_30  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_30 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_31  (
    .i0(inst_dob_i48_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_31 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_32  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_32 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_33  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_33 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_34  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_34 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_35  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_35 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_36  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_36 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_37  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_37 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_38  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_38 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_39  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_39 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_4  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_4 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_40  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_40 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_41  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_41 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_42  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_42 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_43  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_43 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_44  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_44 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_45  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_45 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_46  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_46 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_47  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_47 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_48  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_48 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_49  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_49 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_5  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_5 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_50  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_50 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_51  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_51 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_52  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_52 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_53  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_53 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_54  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_54 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_55  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_55 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_56  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_56 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_57  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_57 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_58  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_58 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_59  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_59 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_6  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_6 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_60  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_60 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_61  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_61 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_62  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_62 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_63  (
    .i0(inst_dob_i64_013),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_63 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_7  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i0_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_7 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_8  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_8 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_9  (
    .i0(inst_dob_i16_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_9 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b13/B0_0 ),
    .i1(\inst_dob_mux_b13/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b13/B0_2 ),
    .i1(\inst_dob_mux_b13/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b13/B0_20 ),
    .i1(\inst_dob_mux_b13/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_10 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b13/B0_22 ),
    .i1(\inst_dob_mux_b13/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_11 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b13/B0_24 ),
    .i1(\inst_dob_mux_b13/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_12 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b13/B0_26 ),
    .i1(\inst_dob_mux_b13/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_13 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b13/B0_28 ),
    .i1(\inst_dob_mux_b13/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_14 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b13/B0_30 ),
    .i1(\inst_dob_mux_b13/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_15 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b13/B0_32 ),
    .i1(\inst_dob_mux_b13/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_16 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b13/B0_34 ),
    .i1(\inst_dob_mux_b13/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_17 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b13/B0_36 ),
    .i1(\inst_dob_mux_b13/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_18 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b13/B0_38 ),
    .i1(\inst_dob_mux_b13/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_19 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b13/B0_4 ),
    .i1(\inst_dob_mux_b13/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_2 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b13/B0_40 ),
    .i1(\inst_dob_mux_b13/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_20 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b13/B0_42 ),
    .i1(\inst_dob_mux_b13/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_21 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b13/B0_44 ),
    .i1(\inst_dob_mux_b13/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_22 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b13/B0_46 ),
    .i1(\inst_dob_mux_b13/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_23 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b13/B0_48 ),
    .i1(\inst_dob_mux_b13/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_24 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b13/B0_50 ),
    .i1(\inst_dob_mux_b13/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_25 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b13/B0_52 ),
    .i1(\inst_dob_mux_b13/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_26 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b13/B0_54 ),
    .i1(\inst_dob_mux_b13/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_27 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b13/B0_56 ),
    .i1(\inst_dob_mux_b13/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_28 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b13/B0_58 ),
    .i1(\inst_dob_mux_b13/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_29 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b13/B0_6 ),
    .i1(\inst_dob_mux_b13/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_3 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b13/B0_60 ),
    .i1(\inst_dob_mux_b13/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_30 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b13/B0_62 ),
    .i1(\inst_dob_mux_b13/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_31 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b13/B0_8 ),
    .i1(\inst_dob_mux_b13/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_4 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b13/B0_10 ),
    .i1(\inst_dob_mux_b13/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_5 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b13/B0_12 ),
    .i1(\inst_dob_mux_b13/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_6 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b13/B0_14 ),
    .i1(\inst_dob_mux_b13/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_7 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b13/B0_16 ),
    .i1(\inst_dob_mux_b13/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_8 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b13/B0_18 ),
    .i1(\inst_dob_mux_b13/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_9 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b13/B1_0 ),
    .i1(\inst_dob_mux_b13/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b13/B1_2 ),
    .i1(\inst_dob_mux_b13/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b13/B1_20 ),
    .i1(\inst_dob_mux_b13/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_10 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b13/B1_22 ),
    .i1(\inst_dob_mux_b13/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_11 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b13/B1_24 ),
    .i1(\inst_dob_mux_b13/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_12 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b13/B1_26 ),
    .i1(\inst_dob_mux_b13/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_13 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b13/B1_28 ),
    .i1(\inst_dob_mux_b13/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_14 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b13/B1_30 ),
    .i1(\inst_dob_mux_b13/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_15 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b13/B1_4 ),
    .i1(\inst_dob_mux_b13/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_2 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b13/B1_6 ),
    .i1(\inst_dob_mux_b13/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_3 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b13/B1_8 ),
    .i1(\inst_dob_mux_b13/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_4 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b13/B1_10 ),
    .i1(\inst_dob_mux_b13/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_5 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b13/B1_12 ),
    .i1(\inst_dob_mux_b13/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_6 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b13/B1_14 ),
    .i1(\inst_dob_mux_b13/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_7 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b13/B1_16 ),
    .i1(\inst_dob_mux_b13/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_8 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b13/B1_18 ),
    .i1(\inst_dob_mux_b13/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b13/B2_9 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b13/B2_0 ),
    .i1(\inst_dob_mux_b13/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b13/B3_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b13/B2_2 ),
    .i1(\inst_dob_mux_b13/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b13/B3_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b13/B2_4 ),
    .i1(\inst_dob_mux_b13/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b13/B3_2 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b13/B2_6 ),
    .i1(\inst_dob_mux_b13/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b13/B3_3 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b13/B2_8 ),
    .i1(\inst_dob_mux_b13/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b13/B3_4 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b13/B2_10 ),
    .i1(\inst_dob_mux_b13/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b13/B3_5 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b13/B2_12 ),
    .i1(\inst_dob_mux_b13/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b13/B3_6 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b13/B2_14 ),
    .i1(\inst_dob_mux_b13/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b13/B3_7 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b13/B3_0 ),
    .i1(\inst_dob_mux_b13/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b13/B4_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b13/B3_2 ),
    .i1(\inst_dob_mux_b13/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b13/B4_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b13/B3_4 ),
    .i1(\inst_dob_mux_b13/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b13/B4_2 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b13/B3_6 ),
    .i1(\inst_dob_mux_b13/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b13/B4_3 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b13/B4_0 ),
    .i1(\inst_dob_mux_b13/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b13/B5_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b13/B4_2 ),
    .i1(\inst_dob_mux_b13/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b13/B5_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b13/B5_0 ),
    .i1(\inst_dob_mux_b13/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[13]));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_0  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_1  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_10  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_10 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_11  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_11 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_12  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_12 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_13  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_13 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_14  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_14 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_15  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_15 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_16  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_16 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_17  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_17 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_18  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_18 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_19  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_19 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_2  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_2 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_20  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_20 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_21  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_21 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_22  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_22 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_23  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i32_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_23 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_24  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_24 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_25  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_25 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_26  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_26 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_27  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_27 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_28  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_28 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_29  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_29 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_3  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_3 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_30  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_30 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_31  (
    .i0(inst_dob_i48_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_31 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_32  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_32 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_33  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_33 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_34  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_34 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_35  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_35 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_36  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_36 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_37  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_37 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_38  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_38 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_39  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_39 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_4  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_4 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_40  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_40 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_41  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_41 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_42  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_42 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_43  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_43 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_44  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_44 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_45  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_45 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_46  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_46 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_47  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_47 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_48  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_48 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_49  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_49 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_5  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_5 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_50  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_50 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_51  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_51 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_52  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_52 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_53  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_53 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_54  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_54 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_55  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_55 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_56  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_56 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_57  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_57 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_58  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_58 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_59  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_59 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_6  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_6 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_60  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_60 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_61  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_61 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_62  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_62 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_63  (
    .i0(inst_dob_i64_014),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_63 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_7  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i0_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_7 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_8  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_8 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_9  (
    .i0(inst_dob_i16_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_9 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b14/B0_0 ),
    .i1(\inst_dob_mux_b14/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b14/B0_2 ),
    .i1(\inst_dob_mux_b14/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b14/B0_20 ),
    .i1(\inst_dob_mux_b14/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_10 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b14/B0_22 ),
    .i1(\inst_dob_mux_b14/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_11 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b14/B0_24 ),
    .i1(\inst_dob_mux_b14/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_12 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b14/B0_26 ),
    .i1(\inst_dob_mux_b14/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_13 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b14/B0_28 ),
    .i1(\inst_dob_mux_b14/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_14 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b14/B0_30 ),
    .i1(\inst_dob_mux_b14/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_15 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b14/B0_32 ),
    .i1(\inst_dob_mux_b14/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_16 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b14/B0_34 ),
    .i1(\inst_dob_mux_b14/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_17 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b14/B0_36 ),
    .i1(\inst_dob_mux_b14/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_18 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b14/B0_38 ),
    .i1(\inst_dob_mux_b14/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_19 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b14/B0_4 ),
    .i1(\inst_dob_mux_b14/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_2 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b14/B0_40 ),
    .i1(\inst_dob_mux_b14/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_20 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b14/B0_42 ),
    .i1(\inst_dob_mux_b14/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_21 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b14/B0_44 ),
    .i1(\inst_dob_mux_b14/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_22 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b14/B0_46 ),
    .i1(\inst_dob_mux_b14/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_23 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b14/B0_48 ),
    .i1(\inst_dob_mux_b14/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_24 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b14/B0_50 ),
    .i1(\inst_dob_mux_b14/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_25 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b14/B0_52 ),
    .i1(\inst_dob_mux_b14/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_26 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b14/B0_54 ),
    .i1(\inst_dob_mux_b14/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_27 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b14/B0_56 ),
    .i1(\inst_dob_mux_b14/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_28 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b14/B0_58 ),
    .i1(\inst_dob_mux_b14/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_29 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b14/B0_6 ),
    .i1(\inst_dob_mux_b14/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_3 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b14/B0_60 ),
    .i1(\inst_dob_mux_b14/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_30 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b14/B0_62 ),
    .i1(\inst_dob_mux_b14/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_31 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b14/B0_8 ),
    .i1(\inst_dob_mux_b14/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_4 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b14/B0_10 ),
    .i1(\inst_dob_mux_b14/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_5 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b14/B0_12 ),
    .i1(\inst_dob_mux_b14/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_6 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b14/B0_14 ),
    .i1(\inst_dob_mux_b14/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_7 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b14/B0_16 ),
    .i1(\inst_dob_mux_b14/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_8 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b14/B0_18 ),
    .i1(\inst_dob_mux_b14/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_9 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b14/B1_0 ),
    .i1(\inst_dob_mux_b14/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b14/B1_2 ),
    .i1(\inst_dob_mux_b14/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b14/B1_20 ),
    .i1(\inst_dob_mux_b14/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_10 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b14/B1_22 ),
    .i1(\inst_dob_mux_b14/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_11 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b14/B1_24 ),
    .i1(\inst_dob_mux_b14/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_12 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b14/B1_26 ),
    .i1(\inst_dob_mux_b14/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_13 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b14/B1_28 ),
    .i1(\inst_dob_mux_b14/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_14 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b14/B1_30 ),
    .i1(\inst_dob_mux_b14/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_15 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b14/B1_4 ),
    .i1(\inst_dob_mux_b14/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_2 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b14/B1_6 ),
    .i1(\inst_dob_mux_b14/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_3 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b14/B1_8 ),
    .i1(\inst_dob_mux_b14/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_4 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b14/B1_10 ),
    .i1(\inst_dob_mux_b14/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_5 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b14/B1_12 ),
    .i1(\inst_dob_mux_b14/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_6 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b14/B1_14 ),
    .i1(\inst_dob_mux_b14/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_7 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b14/B1_16 ),
    .i1(\inst_dob_mux_b14/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_8 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b14/B1_18 ),
    .i1(\inst_dob_mux_b14/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b14/B2_9 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b14/B2_0 ),
    .i1(\inst_dob_mux_b14/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b14/B3_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b14/B2_2 ),
    .i1(\inst_dob_mux_b14/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b14/B3_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b14/B2_4 ),
    .i1(\inst_dob_mux_b14/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b14/B3_2 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b14/B2_6 ),
    .i1(\inst_dob_mux_b14/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b14/B3_3 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b14/B2_8 ),
    .i1(\inst_dob_mux_b14/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b14/B3_4 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b14/B2_10 ),
    .i1(\inst_dob_mux_b14/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b14/B3_5 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b14/B2_12 ),
    .i1(\inst_dob_mux_b14/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b14/B3_6 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b14/B2_14 ),
    .i1(\inst_dob_mux_b14/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b14/B3_7 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b14/B3_0 ),
    .i1(\inst_dob_mux_b14/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b14/B4_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b14/B3_2 ),
    .i1(\inst_dob_mux_b14/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b14/B4_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b14/B3_4 ),
    .i1(\inst_dob_mux_b14/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b14/B4_2 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b14/B3_6 ),
    .i1(\inst_dob_mux_b14/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b14/B4_3 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b14/B4_0 ),
    .i1(\inst_dob_mux_b14/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b14/B5_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b14/B4_2 ),
    .i1(\inst_dob_mux_b14/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b14/B5_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b14/B5_0 ),
    .i1(\inst_dob_mux_b14/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[14]));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_0  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_1  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_10  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_10 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_11  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_11 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_12  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_12 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_13  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_13 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_14  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_14 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_15  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_15 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_16  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_16 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_17  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_17 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_18  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_18 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_19  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_19 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_2  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_2 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_20  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_20 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_21  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_21 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_22  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_22 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_23  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i32_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_23 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_24  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_24 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_25  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_25 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_26  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_26 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_27  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_27 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_28  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_28 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_29  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_29 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_3  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_3 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_30  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_30 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_31  (
    .i0(inst_dob_i48_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_31 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_32  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_32 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_33  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_33 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_34  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_34 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_35  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_35 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_36  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_36 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_37  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_37 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_38  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_38 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_39  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_39 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_4  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_4 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_40  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_40 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_41  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_41 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_42  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_42 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_43  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_43 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_44  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_44 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_45  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_45 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_46  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_46 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_47  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_47 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_48  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_48 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_49  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_49 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_5  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_5 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_50  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_50 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_51  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_51 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_52  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_52 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_53  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_53 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_54  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_54 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_55  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_55 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_56  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_56 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_57  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_57 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_58  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_58 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_59  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_59 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_6  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_6 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_60  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_60 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_61  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_61 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_62  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_62 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_63  (
    .i0(inst_dob_i64_015),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_63 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_7  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i0_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_7 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_8  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_8 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_9  (
    .i0(inst_dob_i16_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_9 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b15/B0_0 ),
    .i1(\inst_dob_mux_b15/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b15/B0_2 ),
    .i1(\inst_dob_mux_b15/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b15/B0_20 ),
    .i1(\inst_dob_mux_b15/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_10 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b15/B0_22 ),
    .i1(\inst_dob_mux_b15/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_11 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b15/B0_24 ),
    .i1(\inst_dob_mux_b15/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_12 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b15/B0_26 ),
    .i1(\inst_dob_mux_b15/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_13 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b15/B0_28 ),
    .i1(\inst_dob_mux_b15/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_14 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b15/B0_30 ),
    .i1(\inst_dob_mux_b15/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_15 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b15/B0_32 ),
    .i1(\inst_dob_mux_b15/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_16 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b15/B0_34 ),
    .i1(\inst_dob_mux_b15/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_17 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b15/B0_36 ),
    .i1(\inst_dob_mux_b15/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_18 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b15/B0_38 ),
    .i1(\inst_dob_mux_b15/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_19 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b15/B0_4 ),
    .i1(\inst_dob_mux_b15/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_2 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b15/B0_40 ),
    .i1(\inst_dob_mux_b15/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_20 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b15/B0_42 ),
    .i1(\inst_dob_mux_b15/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_21 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b15/B0_44 ),
    .i1(\inst_dob_mux_b15/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_22 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b15/B0_46 ),
    .i1(\inst_dob_mux_b15/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_23 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b15/B0_48 ),
    .i1(\inst_dob_mux_b15/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_24 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b15/B0_50 ),
    .i1(\inst_dob_mux_b15/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_25 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b15/B0_52 ),
    .i1(\inst_dob_mux_b15/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_26 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b15/B0_54 ),
    .i1(\inst_dob_mux_b15/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_27 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b15/B0_56 ),
    .i1(\inst_dob_mux_b15/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_28 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b15/B0_58 ),
    .i1(\inst_dob_mux_b15/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_29 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b15/B0_6 ),
    .i1(\inst_dob_mux_b15/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_3 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b15/B0_60 ),
    .i1(\inst_dob_mux_b15/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_30 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b15/B0_62 ),
    .i1(\inst_dob_mux_b15/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_31 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b15/B0_8 ),
    .i1(\inst_dob_mux_b15/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_4 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b15/B0_10 ),
    .i1(\inst_dob_mux_b15/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_5 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b15/B0_12 ),
    .i1(\inst_dob_mux_b15/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_6 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b15/B0_14 ),
    .i1(\inst_dob_mux_b15/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_7 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b15/B0_16 ),
    .i1(\inst_dob_mux_b15/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_8 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b15/B0_18 ),
    .i1(\inst_dob_mux_b15/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_9 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b15/B1_0 ),
    .i1(\inst_dob_mux_b15/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b15/B1_2 ),
    .i1(\inst_dob_mux_b15/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b15/B1_20 ),
    .i1(\inst_dob_mux_b15/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_10 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b15/B1_22 ),
    .i1(\inst_dob_mux_b15/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_11 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b15/B1_24 ),
    .i1(\inst_dob_mux_b15/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_12 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b15/B1_26 ),
    .i1(\inst_dob_mux_b15/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_13 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b15/B1_28 ),
    .i1(\inst_dob_mux_b15/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_14 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b15/B1_30 ),
    .i1(\inst_dob_mux_b15/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_15 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b15/B1_4 ),
    .i1(\inst_dob_mux_b15/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_2 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b15/B1_6 ),
    .i1(\inst_dob_mux_b15/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_3 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b15/B1_8 ),
    .i1(\inst_dob_mux_b15/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_4 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b15/B1_10 ),
    .i1(\inst_dob_mux_b15/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_5 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b15/B1_12 ),
    .i1(\inst_dob_mux_b15/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_6 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b15/B1_14 ),
    .i1(\inst_dob_mux_b15/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_7 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b15/B1_16 ),
    .i1(\inst_dob_mux_b15/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_8 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b15/B1_18 ),
    .i1(\inst_dob_mux_b15/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b15/B2_9 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b15/B2_0 ),
    .i1(\inst_dob_mux_b15/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b15/B3_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b15/B2_2 ),
    .i1(\inst_dob_mux_b15/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b15/B3_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b15/B2_4 ),
    .i1(\inst_dob_mux_b15/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b15/B3_2 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b15/B2_6 ),
    .i1(\inst_dob_mux_b15/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b15/B3_3 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b15/B2_8 ),
    .i1(\inst_dob_mux_b15/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b15/B3_4 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b15/B2_10 ),
    .i1(\inst_dob_mux_b15/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b15/B3_5 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b15/B2_12 ),
    .i1(\inst_dob_mux_b15/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b15/B3_6 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b15/B2_14 ),
    .i1(\inst_dob_mux_b15/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b15/B3_7 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b15/B3_0 ),
    .i1(\inst_dob_mux_b15/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b15/B4_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b15/B3_2 ),
    .i1(\inst_dob_mux_b15/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b15/B4_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b15/B3_4 ),
    .i1(\inst_dob_mux_b15/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b15/B4_2 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b15/B3_6 ),
    .i1(\inst_dob_mux_b15/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b15/B4_3 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b15/B4_0 ),
    .i1(\inst_dob_mux_b15/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b15/B5_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b15/B4_2 ),
    .i1(\inst_dob_mux_b15/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b15/B5_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b15/B5_0 ),
    .i1(\inst_dob_mux_b15/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[15]));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_0  (
    .i0(inst_dob_i0_002),
    .i1(inst_dob_i0_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_1  (
    .i0(inst_dob_i2_002),
    .i1(inst_dob_i2_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_10  (
    .i0(inst_dob_i20_002),
    .i1(inst_dob_i20_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_10 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_11  (
    .i0(inst_dob_i22_002),
    .i1(inst_dob_i22_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_11 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_12  (
    .i0(inst_dob_i24_002),
    .i1(inst_dob_i24_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_12 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_13  (
    .i0(inst_dob_i26_002),
    .i1(inst_dob_i26_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_13 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_14  (
    .i0(inst_dob_i28_002),
    .i1(inst_dob_i28_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_14 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_15  (
    .i0(inst_dob_i30_002),
    .i1(inst_dob_i30_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_15 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_16  (
    .i0(inst_dob_i32_002),
    .i1(inst_dob_i32_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_16 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_17  (
    .i0(inst_dob_i34_002),
    .i1(inst_dob_i34_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_17 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_18  (
    .i0(inst_dob_i36_002),
    .i1(inst_dob_i36_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_18 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_19  (
    .i0(inst_dob_i38_002),
    .i1(inst_dob_i38_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_19 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_2  (
    .i0(inst_dob_i4_002),
    .i1(inst_dob_i4_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_20  (
    .i0(inst_dob_i40_002),
    .i1(inst_dob_i40_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_20 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_21  (
    .i0(inst_dob_i42_002),
    .i1(inst_dob_i42_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_21 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_22  (
    .i0(inst_dob_i44_002),
    .i1(inst_dob_i44_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_22 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_23  (
    .i0(inst_dob_i46_002),
    .i1(inst_dob_i46_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_23 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_24  (
    .i0(inst_dob_i48_002),
    .i1(inst_dob_i48_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_24 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_25  (
    .i0(inst_dob_i50_002),
    .i1(inst_dob_i50_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_25 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_26  (
    .i0(inst_dob_i52_002),
    .i1(inst_dob_i52_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_26 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_27  (
    .i0(inst_dob_i54_002),
    .i1(inst_dob_i54_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_27 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_28  (
    .i0(inst_dob_i56_002),
    .i1(inst_dob_i56_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_28 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_29  (
    .i0(inst_dob_i58_002),
    .i1(inst_dob_i58_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_29 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_3  (
    .i0(inst_dob_i6_002),
    .i1(inst_dob_i6_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_30  (
    .i0(inst_dob_i60_002),
    .i1(inst_dob_i60_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_30 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_31  (
    .i0(inst_dob_i62_002),
    .i1(inst_dob_i62_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_31 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_32  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_32 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_33  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_33 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_34  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_34 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_35  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_35 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_36  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_36 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_37  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_37 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_38  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_38 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_39  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_39 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_4  (
    .i0(inst_dob_i8_002),
    .i1(inst_dob_i8_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_4 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_40  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_40 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_41  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_41 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_42  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_42 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_43  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_43 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_44  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_44 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_45  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_45 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_46  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_46 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_47  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_47 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_48  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_48 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_49  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_49 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_5  (
    .i0(inst_dob_i10_002),
    .i1(inst_dob_i10_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_5 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_50  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_50 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_51  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_51 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_52  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_52 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_53  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_53 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_54  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_54 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_55  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_55 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_56  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_56 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_57  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_57 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_58  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_58 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_59  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_59 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_6  (
    .i0(inst_dob_i12_002),
    .i1(inst_dob_i12_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_6 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_60  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_60 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_61  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_61 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_62  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_62 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_63  (
    .i0(inst_dob_i64_002),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_63 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_7  (
    .i0(inst_dob_i14_002),
    .i1(inst_dob_i14_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_7 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_8  (
    .i0(inst_dob_i16_002),
    .i1(inst_dob_i16_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_8 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_9  (
    .i0(inst_dob_i18_002),
    .i1(inst_dob_i18_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_9 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b2/B0_0 ),
    .i1(\inst_dob_mux_b2/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b2/B0_2 ),
    .i1(\inst_dob_mux_b2/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b2/B0_20 ),
    .i1(\inst_dob_mux_b2/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_10 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b2/B0_22 ),
    .i1(\inst_dob_mux_b2/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_11 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b2/B0_24 ),
    .i1(\inst_dob_mux_b2/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_12 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b2/B0_26 ),
    .i1(\inst_dob_mux_b2/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_13 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b2/B0_28 ),
    .i1(\inst_dob_mux_b2/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_14 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b2/B0_30 ),
    .i1(\inst_dob_mux_b2/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_15 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b2/B0_32 ),
    .i1(\inst_dob_mux_b2/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_16 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b2/B0_34 ),
    .i1(\inst_dob_mux_b2/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_17 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b2/B0_36 ),
    .i1(\inst_dob_mux_b2/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_18 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b2/B0_38 ),
    .i1(\inst_dob_mux_b2/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_19 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b2/B0_4 ),
    .i1(\inst_dob_mux_b2/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b2/B0_40 ),
    .i1(\inst_dob_mux_b2/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_20 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b2/B0_42 ),
    .i1(\inst_dob_mux_b2/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_21 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b2/B0_44 ),
    .i1(\inst_dob_mux_b2/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_22 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b2/B0_46 ),
    .i1(\inst_dob_mux_b2/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_23 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b2/B0_48 ),
    .i1(\inst_dob_mux_b2/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_24 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b2/B0_50 ),
    .i1(\inst_dob_mux_b2/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_25 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b2/B0_52 ),
    .i1(\inst_dob_mux_b2/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_26 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b2/B0_54 ),
    .i1(\inst_dob_mux_b2/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_27 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b2/B0_56 ),
    .i1(\inst_dob_mux_b2/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_28 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b2/B0_58 ),
    .i1(\inst_dob_mux_b2/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_29 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b2/B0_6 ),
    .i1(\inst_dob_mux_b2/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b2/B0_60 ),
    .i1(\inst_dob_mux_b2/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_30 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b2/B0_62 ),
    .i1(\inst_dob_mux_b2/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_31 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b2/B0_8 ),
    .i1(\inst_dob_mux_b2/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_4 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b2/B0_10 ),
    .i1(\inst_dob_mux_b2/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_5 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b2/B0_12 ),
    .i1(\inst_dob_mux_b2/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_6 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b2/B0_14 ),
    .i1(\inst_dob_mux_b2/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_7 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b2/B0_16 ),
    .i1(\inst_dob_mux_b2/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_8 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b2/B0_18 ),
    .i1(\inst_dob_mux_b2/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_9 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b2/B1_0 ),
    .i1(\inst_dob_mux_b2/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b2/B1_2 ),
    .i1(\inst_dob_mux_b2/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b2/B1_20 ),
    .i1(\inst_dob_mux_b2/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_10 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b2/B1_22 ),
    .i1(\inst_dob_mux_b2/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_11 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b2/B1_24 ),
    .i1(\inst_dob_mux_b2/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_12 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b2/B1_26 ),
    .i1(\inst_dob_mux_b2/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_13 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b2/B1_28 ),
    .i1(\inst_dob_mux_b2/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_14 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b2/B1_30 ),
    .i1(\inst_dob_mux_b2/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_15 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b2/B1_4 ),
    .i1(\inst_dob_mux_b2/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b2/B1_6 ),
    .i1(\inst_dob_mux_b2/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b2/B1_8 ),
    .i1(\inst_dob_mux_b2/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_4 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b2/B1_10 ),
    .i1(\inst_dob_mux_b2/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_5 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b2/B1_12 ),
    .i1(\inst_dob_mux_b2/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_6 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b2/B1_14 ),
    .i1(\inst_dob_mux_b2/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_7 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b2/B1_16 ),
    .i1(\inst_dob_mux_b2/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_8 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b2/B1_18 ),
    .i1(\inst_dob_mux_b2/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_9 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b2/B2_0 ),
    .i1(\inst_dob_mux_b2/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b2/B3_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b2/B2_2 ),
    .i1(\inst_dob_mux_b2/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b2/B3_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b2/B2_4 ),
    .i1(\inst_dob_mux_b2/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b2/B3_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b2/B2_6 ),
    .i1(\inst_dob_mux_b2/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b2/B3_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b2/B2_8 ),
    .i1(\inst_dob_mux_b2/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b2/B3_4 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b2/B2_10 ),
    .i1(\inst_dob_mux_b2/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b2/B3_5 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b2/B2_12 ),
    .i1(\inst_dob_mux_b2/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b2/B3_6 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b2/B2_14 ),
    .i1(\inst_dob_mux_b2/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b2/B3_7 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b2/B3_0 ),
    .i1(\inst_dob_mux_b2/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b2/B4_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b2/B3_2 ),
    .i1(\inst_dob_mux_b2/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b2/B4_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b2/B3_4 ),
    .i1(\inst_dob_mux_b2/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b2/B4_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b2/B3_6 ),
    .i1(\inst_dob_mux_b2/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b2/B4_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b2/B4_0 ),
    .i1(\inst_dob_mux_b2/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b2/B5_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b2/B4_2 ),
    .i1(\inst_dob_mux_b2/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b2/B5_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b2/B5_0 ),
    .i1(\inst_dob_mux_b2/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[2]));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_0  (
    .i0(inst_dob_i0_003),
    .i1(inst_dob_i0_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_1  (
    .i0(inst_dob_i2_003),
    .i1(inst_dob_i2_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_10  (
    .i0(inst_dob_i20_003),
    .i1(inst_dob_i20_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_10 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_11  (
    .i0(inst_dob_i22_003),
    .i1(inst_dob_i22_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_11 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_12  (
    .i0(inst_dob_i24_003),
    .i1(inst_dob_i24_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_12 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_13  (
    .i0(inst_dob_i26_003),
    .i1(inst_dob_i26_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_13 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_14  (
    .i0(inst_dob_i28_003),
    .i1(inst_dob_i28_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_14 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_15  (
    .i0(inst_dob_i30_003),
    .i1(inst_dob_i30_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_15 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_16  (
    .i0(inst_dob_i32_003),
    .i1(inst_dob_i32_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_16 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_17  (
    .i0(inst_dob_i34_003),
    .i1(inst_dob_i34_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_17 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_18  (
    .i0(inst_dob_i36_003),
    .i1(inst_dob_i36_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_18 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_19  (
    .i0(inst_dob_i38_003),
    .i1(inst_dob_i38_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_19 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_2  (
    .i0(inst_dob_i4_003),
    .i1(inst_dob_i4_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_20  (
    .i0(inst_dob_i40_003),
    .i1(inst_dob_i40_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_20 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_21  (
    .i0(inst_dob_i42_003),
    .i1(inst_dob_i42_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_21 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_22  (
    .i0(inst_dob_i44_003),
    .i1(inst_dob_i44_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_22 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_23  (
    .i0(inst_dob_i46_003),
    .i1(inst_dob_i46_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_23 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_24  (
    .i0(inst_dob_i48_003),
    .i1(inst_dob_i48_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_24 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_25  (
    .i0(inst_dob_i50_003),
    .i1(inst_dob_i50_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_25 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_26  (
    .i0(inst_dob_i52_003),
    .i1(inst_dob_i52_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_26 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_27  (
    .i0(inst_dob_i54_003),
    .i1(inst_dob_i54_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_27 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_28  (
    .i0(inst_dob_i56_003),
    .i1(inst_dob_i56_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_28 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_29  (
    .i0(inst_dob_i58_003),
    .i1(inst_dob_i58_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_29 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_3  (
    .i0(inst_dob_i6_003),
    .i1(inst_dob_i6_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_30  (
    .i0(inst_dob_i60_003),
    .i1(inst_dob_i60_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_30 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_31  (
    .i0(inst_dob_i62_003),
    .i1(inst_dob_i62_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_31 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_32  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_32 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_33  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_33 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_34  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_34 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_35  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_35 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_36  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_36 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_37  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_37 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_38  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_38 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_39  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_39 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_4  (
    .i0(inst_dob_i8_003),
    .i1(inst_dob_i8_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_4 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_40  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_40 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_41  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_41 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_42  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_42 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_43  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_43 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_44  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_44 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_45  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_45 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_46  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_46 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_47  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_47 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_48  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_48 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_49  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_49 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_5  (
    .i0(inst_dob_i10_003),
    .i1(inst_dob_i10_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_5 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_50  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_50 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_51  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_51 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_52  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_52 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_53  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_53 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_54  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_54 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_55  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_55 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_56  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_56 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_57  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_57 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_58  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_58 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_59  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_59 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_6  (
    .i0(inst_dob_i12_003),
    .i1(inst_dob_i12_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_6 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_60  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_60 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_61  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_61 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_62  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_62 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_63  (
    .i0(inst_dob_i64_003),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_63 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_7  (
    .i0(inst_dob_i14_003),
    .i1(inst_dob_i14_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_7 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_8  (
    .i0(inst_dob_i16_003),
    .i1(inst_dob_i16_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_8 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_9  (
    .i0(inst_dob_i18_003),
    .i1(inst_dob_i18_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_9 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b3/B0_0 ),
    .i1(\inst_dob_mux_b3/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b3/B0_2 ),
    .i1(\inst_dob_mux_b3/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b3/B0_20 ),
    .i1(\inst_dob_mux_b3/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_10 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b3/B0_22 ),
    .i1(\inst_dob_mux_b3/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_11 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b3/B0_24 ),
    .i1(\inst_dob_mux_b3/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_12 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b3/B0_26 ),
    .i1(\inst_dob_mux_b3/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_13 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b3/B0_28 ),
    .i1(\inst_dob_mux_b3/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_14 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b3/B0_30 ),
    .i1(\inst_dob_mux_b3/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_15 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b3/B0_32 ),
    .i1(\inst_dob_mux_b3/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_16 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b3/B0_34 ),
    .i1(\inst_dob_mux_b3/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_17 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b3/B0_36 ),
    .i1(\inst_dob_mux_b3/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_18 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b3/B0_38 ),
    .i1(\inst_dob_mux_b3/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_19 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b3/B0_4 ),
    .i1(\inst_dob_mux_b3/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b3/B0_40 ),
    .i1(\inst_dob_mux_b3/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_20 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b3/B0_42 ),
    .i1(\inst_dob_mux_b3/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_21 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b3/B0_44 ),
    .i1(\inst_dob_mux_b3/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_22 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b3/B0_46 ),
    .i1(\inst_dob_mux_b3/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_23 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b3/B0_48 ),
    .i1(\inst_dob_mux_b3/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_24 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b3/B0_50 ),
    .i1(\inst_dob_mux_b3/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_25 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b3/B0_52 ),
    .i1(\inst_dob_mux_b3/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_26 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b3/B0_54 ),
    .i1(\inst_dob_mux_b3/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_27 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b3/B0_56 ),
    .i1(\inst_dob_mux_b3/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_28 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b3/B0_58 ),
    .i1(\inst_dob_mux_b3/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_29 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b3/B0_6 ),
    .i1(\inst_dob_mux_b3/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b3/B0_60 ),
    .i1(\inst_dob_mux_b3/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_30 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b3/B0_62 ),
    .i1(\inst_dob_mux_b3/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_31 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b3/B0_8 ),
    .i1(\inst_dob_mux_b3/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_4 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b3/B0_10 ),
    .i1(\inst_dob_mux_b3/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_5 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b3/B0_12 ),
    .i1(\inst_dob_mux_b3/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_6 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b3/B0_14 ),
    .i1(\inst_dob_mux_b3/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_7 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b3/B0_16 ),
    .i1(\inst_dob_mux_b3/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_8 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b3/B0_18 ),
    .i1(\inst_dob_mux_b3/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_9 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b3/B1_0 ),
    .i1(\inst_dob_mux_b3/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b3/B1_2 ),
    .i1(\inst_dob_mux_b3/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b3/B1_20 ),
    .i1(\inst_dob_mux_b3/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_10 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b3/B1_22 ),
    .i1(\inst_dob_mux_b3/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_11 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b3/B1_24 ),
    .i1(\inst_dob_mux_b3/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_12 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b3/B1_26 ),
    .i1(\inst_dob_mux_b3/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_13 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b3/B1_28 ),
    .i1(\inst_dob_mux_b3/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_14 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b3/B1_30 ),
    .i1(\inst_dob_mux_b3/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_15 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b3/B1_4 ),
    .i1(\inst_dob_mux_b3/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b3/B1_6 ),
    .i1(\inst_dob_mux_b3/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b3/B1_8 ),
    .i1(\inst_dob_mux_b3/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_4 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b3/B1_10 ),
    .i1(\inst_dob_mux_b3/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_5 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b3/B1_12 ),
    .i1(\inst_dob_mux_b3/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_6 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b3/B1_14 ),
    .i1(\inst_dob_mux_b3/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_7 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b3/B1_16 ),
    .i1(\inst_dob_mux_b3/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_8 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b3/B1_18 ),
    .i1(\inst_dob_mux_b3/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_9 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b3/B2_0 ),
    .i1(\inst_dob_mux_b3/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b3/B3_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b3/B2_2 ),
    .i1(\inst_dob_mux_b3/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b3/B3_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b3/B2_4 ),
    .i1(\inst_dob_mux_b3/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b3/B3_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b3/B2_6 ),
    .i1(\inst_dob_mux_b3/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b3/B3_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b3/B2_8 ),
    .i1(\inst_dob_mux_b3/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b3/B3_4 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b3/B2_10 ),
    .i1(\inst_dob_mux_b3/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b3/B3_5 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b3/B2_12 ),
    .i1(\inst_dob_mux_b3/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b3/B3_6 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b3/B2_14 ),
    .i1(\inst_dob_mux_b3/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b3/B3_7 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b3/B3_0 ),
    .i1(\inst_dob_mux_b3/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b3/B4_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b3/B3_2 ),
    .i1(\inst_dob_mux_b3/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b3/B4_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b3/B3_4 ),
    .i1(\inst_dob_mux_b3/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b3/B4_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b3/B3_6 ),
    .i1(\inst_dob_mux_b3/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b3/B4_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b3/B4_0 ),
    .i1(\inst_dob_mux_b3/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b3/B5_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b3/B4_2 ),
    .i1(\inst_dob_mux_b3/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b3/B5_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b3/B5_0 ),
    .i1(\inst_dob_mux_b3/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[3]));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_0  (
    .i0(inst_dob_i0_004),
    .i1(inst_dob_i0_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_1  (
    .i0(inst_dob_i2_004),
    .i1(inst_dob_i2_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_10  (
    .i0(inst_dob_i20_004),
    .i1(inst_dob_i20_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_10 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_11  (
    .i0(inst_dob_i22_004),
    .i1(inst_dob_i22_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_11 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_12  (
    .i0(inst_dob_i24_004),
    .i1(inst_dob_i24_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_12 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_13  (
    .i0(inst_dob_i26_004),
    .i1(inst_dob_i26_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_13 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_14  (
    .i0(inst_dob_i28_004),
    .i1(inst_dob_i28_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_14 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_15  (
    .i0(inst_dob_i30_004),
    .i1(inst_dob_i30_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_15 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_16  (
    .i0(inst_dob_i32_004),
    .i1(inst_dob_i32_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_16 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_17  (
    .i0(inst_dob_i34_004),
    .i1(inst_dob_i34_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_17 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_18  (
    .i0(inst_dob_i36_004),
    .i1(inst_dob_i36_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_18 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_19  (
    .i0(inst_dob_i38_004),
    .i1(inst_dob_i38_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_19 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_2  (
    .i0(inst_dob_i4_004),
    .i1(inst_dob_i4_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_20  (
    .i0(inst_dob_i40_004),
    .i1(inst_dob_i40_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_20 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_21  (
    .i0(inst_dob_i42_004),
    .i1(inst_dob_i42_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_21 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_22  (
    .i0(inst_dob_i44_004),
    .i1(inst_dob_i44_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_22 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_23  (
    .i0(inst_dob_i46_004),
    .i1(inst_dob_i46_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_23 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_24  (
    .i0(inst_dob_i48_004),
    .i1(inst_dob_i48_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_24 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_25  (
    .i0(inst_dob_i50_004),
    .i1(inst_dob_i50_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_25 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_26  (
    .i0(inst_dob_i52_004),
    .i1(inst_dob_i52_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_26 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_27  (
    .i0(inst_dob_i54_004),
    .i1(inst_dob_i54_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_27 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_28  (
    .i0(inst_dob_i56_004),
    .i1(inst_dob_i56_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_28 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_29  (
    .i0(inst_dob_i58_004),
    .i1(inst_dob_i58_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_29 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_3  (
    .i0(inst_dob_i6_004),
    .i1(inst_dob_i6_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_30  (
    .i0(inst_dob_i60_004),
    .i1(inst_dob_i60_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_30 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_31  (
    .i0(inst_dob_i62_004),
    .i1(inst_dob_i62_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_31 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_32  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_32 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_33  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_33 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_34  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_34 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_35  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_35 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_36  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_36 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_37  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_37 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_38  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_38 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_39  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_39 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_4  (
    .i0(inst_dob_i8_004),
    .i1(inst_dob_i8_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_4 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_40  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_40 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_41  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_41 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_42  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_42 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_43  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_43 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_44  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_44 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_45  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_45 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_46  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_46 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_47  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_47 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_48  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_48 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_49  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_49 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_5  (
    .i0(inst_dob_i10_004),
    .i1(inst_dob_i10_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_5 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_50  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_50 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_51  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_51 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_52  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_52 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_53  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_53 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_54  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_54 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_55  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_55 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_56  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_56 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_57  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_57 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_58  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_58 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_59  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_59 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_6  (
    .i0(inst_dob_i12_004),
    .i1(inst_dob_i12_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_6 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_60  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_60 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_61  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_61 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_62  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_62 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_63  (
    .i0(inst_dob_i64_004),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_63 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_7  (
    .i0(inst_dob_i14_004),
    .i1(inst_dob_i14_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_7 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_8  (
    .i0(inst_dob_i16_004),
    .i1(inst_dob_i16_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_8 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_9  (
    .i0(inst_dob_i18_004),
    .i1(inst_dob_i18_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_9 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b4/B0_0 ),
    .i1(\inst_dob_mux_b4/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b4/B0_2 ),
    .i1(\inst_dob_mux_b4/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b4/B0_20 ),
    .i1(\inst_dob_mux_b4/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_10 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b4/B0_22 ),
    .i1(\inst_dob_mux_b4/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_11 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b4/B0_24 ),
    .i1(\inst_dob_mux_b4/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_12 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b4/B0_26 ),
    .i1(\inst_dob_mux_b4/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_13 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b4/B0_28 ),
    .i1(\inst_dob_mux_b4/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_14 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b4/B0_30 ),
    .i1(\inst_dob_mux_b4/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_15 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b4/B0_32 ),
    .i1(\inst_dob_mux_b4/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_16 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b4/B0_34 ),
    .i1(\inst_dob_mux_b4/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_17 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b4/B0_36 ),
    .i1(\inst_dob_mux_b4/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_18 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b4/B0_38 ),
    .i1(\inst_dob_mux_b4/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_19 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b4/B0_4 ),
    .i1(\inst_dob_mux_b4/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b4/B0_40 ),
    .i1(\inst_dob_mux_b4/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_20 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b4/B0_42 ),
    .i1(\inst_dob_mux_b4/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_21 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b4/B0_44 ),
    .i1(\inst_dob_mux_b4/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_22 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b4/B0_46 ),
    .i1(\inst_dob_mux_b4/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_23 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b4/B0_48 ),
    .i1(\inst_dob_mux_b4/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_24 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b4/B0_50 ),
    .i1(\inst_dob_mux_b4/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_25 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b4/B0_52 ),
    .i1(\inst_dob_mux_b4/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_26 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b4/B0_54 ),
    .i1(\inst_dob_mux_b4/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_27 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b4/B0_56 ),
    .i1(\inst_dob_mux_b4/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_28 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b4/B0_58 ),
    .i1(\inst_dob_mux_b4/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_29 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b4/B0_6 ),
    .i1(\inst_dob_mux_b4/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b4/B0_60 ),
    .i1(\inst_dob_mux_b4/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_30 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b4/B0_62 ),
    .i1(\inst_dob_mux_b4/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_31 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b4/B0_8 ),
    .i1(\inst_dob_mux_b4/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_4 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b4/B0_10 ),
    .i1(\inst_dob_mux_b4/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_5 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b4/B0_12 ),
    .i1(\inst_dob_mux_b4/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_6 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b4/B0_14 ),
    .i1(\inst_dob_mux_b4/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_7 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b4/B0_16 ),
    .i1(\inst_dob_mux_b4/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_8 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b4/B0_18 ),
    .i1(\inst_dob_mux_b4/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_9 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b4/B1_0 ),
    .i1(\inst_dob_mux_b4/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b4/B1_2 ),
    .i1(\inst_dob_mux_b4/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b4/B1_20 ),
    .i1(\inst_dob_mux_b4/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_10 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b4/B1_22 ),
    .i1(\inst_dob_mux_b4/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_11 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b4/B1_24 ),
    .i1(\inst_dob_mux_b4/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_12 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b4/B1_26 ),
    .i1(\inst_dob_mux_b4/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_13 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b4/B1_28 ),
    .i1(\inst_dob_mux_b4/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_14 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b4/B1_30 ),
    .i1(\inst_dob_mux_b4/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_15 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b4/B1_4 ),
    .i1(\inst_dob_mux_b4/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b4/B1_6 ),
    .i1(\inst_dob_mux_b4/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b4/B1_8 ),
    .i1(\inst_dob_mux_b4/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_4 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b4/B1_10 ),
    .i1(\inst_dob_mux_b4/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_5 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b4/B1_12 ),
    .i1(\inst_dob_mux_b4/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_6 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b4/B1_14 ),
    .i1(\inst_dob_mux_b4/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_7 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b4/B1_16 ),
    .i1(\inst_dob_mux_b4/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_8 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b4/B1_18 ),
    .i1(\inst_dob_mux_b4/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_9 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b4/B2_0 ),
    .i1(\inst_dob_mux_b4/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b4/B3_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b4/B2_2 ),
    .i1(\inst_dob_mux_b4/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b4/B3_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b4/B2_4 ),
    .i1(\inst_dob_mux_b4/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b4/B3_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b4/B2_6 ),
    .i1(\inst_dob_mux_b4/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b4/B3_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b4/B2_8 ),
    .i1(\inst_dob_mux_b4/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b4/B3_4 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b4/B2_10 ),
    .i1(\inst_dob_mux_b4/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b4/B3_5 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b4/B2_12 ),
    .i1(\inst_dob_mux_b4/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b4/B3_6 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b4/B2_14 ),
    .i1(\inst_dob_mux_b4/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b4/B3_7 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b4/B3_0 ),
    .i1(\inst_dob_mux_b4/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b4/B4_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b4/B3_2 ),
    .i1(\inst_dob_mux_b4/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b4/B4_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b4/B3_4 ),
    .i1(\inst_dob_mux_b4/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b4/B4_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b4/B3_6 ),
    .i1(\inst_dob_mux_b4/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b4/B4_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b4/B4_0 ),
    .i1(\inst_dob_mux_b4/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b4/B5_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b4/B4_2 ),
    .i1(\inst_dob_mux_b4/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b4/B5_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b4/B5_0 ),
    .i1(\inst_dob_mux_b4/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[4]));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_0  (
    .i0(inst_dob_i0_005),
    .i1(inst_dob_i0_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_1  (
    .i0(inst_dob_i2_005),
    .i1(inst_dob_i2_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_10  (
    .i0(inst_dob_i20_005),
    .i1(inst_dob_i20_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_10 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_11  (
    .i0(inst_dob_i22_005),
    .i1(inst_dob_i22_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_11 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_12  (
    .i0(inst_dob_i24_005),
    .i1(inst_dob_i24_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_12 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_13  (
    .i0(inst_dob_i26_005),
    .i1(inst_dob_i26_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_13 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_14  (
    .i0(inst_dob_i28_005),
    .i1(inst_dob_i28_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_14 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_15  (
    .i0(inst_dob_i30_005),
    .i1(inst_dob_i30_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_15 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_16  (
    .i0(inst_dob_i32_005),
    .i1(inst_dob_i32_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_16 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_17  (
    .i0(inst_dob_i34_005),
    .i1(inst_dob_i34_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_17 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_18  (
    .i0(inst_dob_i36_005),
    .i1(inst_dob_i36_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_18 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_19  (
    .i0(inst_dob_i38_005),
    .i1(inst_dob_i38_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_19 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_2  (
    .i0(inst_dob_i4_005),
    .i1(inst_dob_i4_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_20  (
    .i0(inst_dob_i40_005),
    .i1(inst_dob_i40_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_20 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_21  (
    .i0(inst_dob_i42_005),
    .i1(inst_dob_i42_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_21 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_22  (
    .i0(inst_dob_i44_005),
    .i1(inst_dob_i44_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_22 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_23  (
    .i0(inst_dob_i46_005),
    .i1(inst_dob_i46_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_23 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_24  (
    .i0(inst_dob_i48_005),
    .i1(inst_dob_i48_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_24 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_25  (
    .i0(inst_dob_i50_005),
    .i1(inst_dob_i50_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_25 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_26  (
    .i0(inst_dob_i52_005),
    .i1(inst_dob_i52_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_26 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_27  (
    .i0(inst_dob_i54_005),
    .i1(inst_dob_i54_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_27 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_28  (
    .i0(inst_dob_i56_005),
    .i1(inst_dob_i56_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_28 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_29  (
    .i0(inst_dob_i58_005),
    .i1(inst_dob_i58_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_29 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_3  (
    .i0(inst_dob_i6_005),
    .i1(inst_dob_i6_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_30  (
    .i0(inst_dob_i60_005),
    .i1(inst_dob_i60_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_30 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_31  (
    .i0(inst_dob_i62_005),
    .i1(inst_dob_i62_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_31 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_32  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_32 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_33  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_33 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_34  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_34 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_35  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_35 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_36  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_36 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_37  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_37 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_38  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_38 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_39  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_39 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_4  (
    .i0(inst_dob_i8_005),
    .i1(inst_dob_i8_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_4 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_40  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_40 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_41  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_41 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_42  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_42 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_43  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_43 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_44  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_44 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_45  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_45 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_46  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_46 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_47  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_47 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_48  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_48 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_49  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_49 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_5  (
    .i0(inst_dob_i10_005),
    .i1(inst_dob_i10_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_5 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_50  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_50 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_51  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_51 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_52  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_52 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_53  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_53 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_54  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_54 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_55  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_55 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_56  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_56 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_57  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_57 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_58  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_58 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_59  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_59 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_6  (
    .i0(inst_dob_i12_005),
    .i1(inst_dob_i12_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_6 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_60  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_60 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_61  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_61 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_62  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_62 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_63  (
    .i0(inst_dob_i64_005),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_63 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_7  (
    .i0(inst_dob_i14_005),
    .i1(inst_dob_i14_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_7 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_8  (
    .i0(inst_dob_i16_005),
    .i1(inst_dob_i16_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_8 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_9  (
    .i0(inst_dob_i18_005),
    .i1(inst_dob_i18_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_9 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b5/B0_0 ),
    .i1(\inst_dob_mux_b5/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b5/B0_2 ),
    .i1(\inst_dob_mux_b5/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b5/B0_20 ),
    .i1(\inst_dob_mux_b5/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_10 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b5/B0_22 ),
    .i1(\inst_dob_mux_b5/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_11 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b5/B0_24 ),
    .i1(\inst_dob_mux_b5/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_12 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b5/B0_26 ),
    .i1(\inst_dob_mux_b5/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_13 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b5/B0_28 ),
    .i1(\inst_dob_mux_b5/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_14 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b5/B0_30 ),
    .i1(\inst_dob_mux_b5/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_15 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b5/B0_32 ),
    .i1(\inst_dob_mux_b5/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_16 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b5/B0_34 ),
    .i1(\inst_dob_mux_b5/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_17 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b5/B0_36 ),
    .i1(\inst_dob_mux_b5/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_18 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b5/B0_38 ),
    .i1(\inst_dob_mux_b5/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_19 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b5/B0_4 ),
    .i1(\inst_dob_mux_b5/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b5/B0_40 ),
    .i1(\inst_dob_mux_b5/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_20 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b5/B0_42 ),
    .i1(\inst_dob_mux_b5/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_21 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b5/B0_44 ),
    .i1(\inst_dob_mux_b5/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_22 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b5/B0_46 ),
    .i1(\inst_dob_mux_b5/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_23 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b5/B0_48 ),
    .i1(\inst_dob_mux_b5/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_24 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b5/B0_50 ),
    .i1(\inst_dob_mux_b5/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_25 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b5/B0_52 ),
    .i1(\inst_dob_mux_b5/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_26 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b5/B0_54 ),
    .i1(\inst_dob_mux_b5/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_27 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b5/B0_56 ),
    .i1(\inst_dob_mux_b5/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_28 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b5/B0_58 ),
    .i1(\inst_dob_mux_b5/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_29 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b5/B0_6 ),
    .i1(\inst_dob_mux_b5/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b5/B0_60 ),
    .i1(\inst_dob_mux_b5/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_30 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b5/B0_62 ),
    .i1(\inst_dob_mux_b5/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_31 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b5/B0_8 ),
    .i1(\inst_dob_mux_b5/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_4 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b5/B0_10 ),
    .i1(\inst_dob_mux_b5/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_5 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b5/B0_12 ),
    .i1(\inst_dob_mux_b5/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_6 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b5/B0_14 ),
    .i1(\inst_dob_mux_b5/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_7 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b5/B0_16 ),
    .i1(\inst_dob_mux_b5/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_8 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b5/B0_18 ),
    .i1(\inst_dob_mux_b5/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_9 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b5/B1_0 ),
    .i1(\inst_dob_mux_b5/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b5/B1_2 ),
    .i1(\inst_dob_mux_b5/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b5/B1_20 ),
    .i1(\inst_dob_mux_b5/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_10 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b5/B1_22 ),
    .i1(\inst_dob_mux_b5/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_11 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b5/B1_24 ),
    .i1(\inst_dob_mux_b5/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_12 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b5/B1_26 ),
    .i1(\inst_dob_mux_b5/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_13 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b5/B1_28 ),
    .i1(\inst_dob_mux_b5/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_14 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b5/B1_30 ),
    .i1(\inst_dob_mux_b5/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_15 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b5/B1_4 ),
    .i1(\inst_dob_mux_b5/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b5/B1_6 ),
    .i1(\inst_dob_mux_b5/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b5/B1_8 ),
    .i1(\inst_dob_mux_b5/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_4 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b5/B1_10 ),
    .i1(\inst_dob_mux_b5/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_5 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b5/B1_12 ),
    .i1(\inst_dob_mux_b5/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_6 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b5/B1_14 ),
    .i1(\inst_dob_mux_b5/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_7 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b5/B1_16 ),
    .i1(\inst_dob_mux_b5/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_8 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b5/B1_18 ),
    .i1(\inst_dob_mux_b5/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_9 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b5/B2_0 ),
    .i1(\inst_dob_mux_b5/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b5/B3_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b5/B2_2 ),
    .i1(\inst_dob_mux_b5/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b5/B3_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b5/B2_4 ),
    .i1(\inst_dob_mux_b5/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b5/B3_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b5/B2_6 ),
    .i1(\inst_dob_mux_b5/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b5/B3_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b5/B2_8 ),
    .i1(\inst_dob_mux_b5/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b5/B3_4 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b5/B2_10 ),
    .i1(\inst_dob_mux_b5/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b5/B3_5 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b5/B2_12 ),
    .i1(\inst_dob_mux_b5/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b5/B3_6 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b5/B2_14 ),
    .i1(\inst_dob_mux_b5/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b5/B3_7 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b5/B3_0 ),
    .i1(\inst_dob_mux_b5/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b5/B4_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b5/B3_2 ),
    .i1(\inst_dob_mux_b5/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b5/B4_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b5/B3_4 ),
    .i1(\inst_dob_mux_b5/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b5/B4_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b5/B3_6 ),
    .i1(\inst_dob_mux_b5/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b5/B4_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b5/B4_0 ),
    .i1(\inst_dob_mux_b5/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b5/B5_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b5/B4_2 ),
    .i1(\inst_dob_mux_b5/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b5/B5_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b5/B5_0 ),
    .i1(\inst_dob_mux_b5/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[5]));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_0  (
    .i0(inst_dob_i0_006),
    .i1(inst_dob_i0_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_1  (
    .i0(inst_dob_i2_006),
    .i1(inst_dob_i2_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_10  (
    .i0(inst_dob_i20_006),
    .i1(inst_dob_i20_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_10 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_11  (
    .i0(inst_dob_i22_006),
    .i1(inst_dob_i22_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_11 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_12  (
    .i0(inst_dob_i24_006),
    .i1(inst_dob_i24_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_12 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_13  (
    .i0(inst_dob_i26_006),
    .i1(inst_dob_i26_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_13 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_14  (
    .i0(inst_dob_i28_006),
    .i1(inst_dob_i28_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_14 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_15  (
    .i0(inst_dob_i30_006),
    .i1(inst_dob_i30_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_15 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_16  (
    .i0(inst_dob_i32_006),
    .i1(inst_dob_i32_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_16 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_17  (
    .i0(inst_dob_i34_006),
    .i1(inst_dob_i34_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_17 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_18  (
    .i0(inst_dob_i36_006),
    .i1(inst_dob_i36_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_18 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_19  (
    .i0(inst_dob_i38_006),
    .i1(inst_dob_i38_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_19 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_2  (
    .i0(inst_dob_i4_006),
    .i1(inst_dob_i4_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_20  (
    .i0(inst_dob_i40_006),
    .i1(inst_dob_i40_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_20 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_21  (
    .i0(inst_dob_i42_006),
    .i1(inst_dob_i42_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_21 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_22  (
    .i0(inst_dob_i44_006),
    .i1(inst_dob_i44_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_22 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_23  (
    .i0(inst_dob_i46_006),
    .i1(inst_dob_i46_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_23 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_24  (
    .i0(inst_dob_i48_006),
    .i1(inst_dob_i48_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_24 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_25  (
    .i0(inst_dob_i50_006),
    .i1(inst_dob_i50_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_25 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_26  (
    .i0(inst_dob_i52_006),
    .i1(inst_dob_i52_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_26 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_27  (
    .i0(inst_dob_i54_006),
    .i1(inst_dob_i54_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_27 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_28  (
    .i0(inst_dob_i56_006),
    .i1(inst_dob_i56_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_28 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_29  (
    .i0(inst_dob_i58_006),
    .i1(inst_dob_i58_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_29 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_3  (
    .i0(inst_dob_i6_006),
    .i1(inst_dob_i6_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_30  (
    .i0(inst_dob_i60_006),
    .i1(inst_dob_i60_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_30 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_31  (
    .i0(inst_dob_i62_006),
    .i1(inst_dob_i62_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_31 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_32  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_32 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_33  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_33 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_34  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_34 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_35  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_35 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_36  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_36 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_37  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_37 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_38  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_38 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_39  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_39 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_4  (
    .i0(inst_dob_i8_006),
    .i1(inst_dob_i8_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_4 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_40  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_40 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_41  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_41 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_42  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_42 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_43  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_43 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_44  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_44 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_45  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_45 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_46  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_46 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_47  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_47 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_48  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_48 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_49  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_49 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_5  (
    .i0(inst_dob_i10_006),
    .i1(inst_dob_i10_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_5 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_50  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_50 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_51  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_51 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_52  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_52 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_53  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_53 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_54  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_54 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_55  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_55 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_56  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_56 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_57  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_57 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_58  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_58 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_59  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_59 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_6  (
    .i0(inst_dob_i12_006),
    .i1(inst_dob_i12_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_6 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_60  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_60 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_61  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_61 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_62  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_62 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_63  (
    .i0(inst_dob_i64_006),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_63 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_7  (
    .i0(inst_dob_i14_006),
    .i1(inst_dob_i14_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_7 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_8  (
    .i0(inst_dob_i16_006),
    .i1(inst_dob_i16_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_8 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_9  (
    .i0(inst_dob_i18_006),
    .i1(inst_dob_i18_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_9 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b6/B0_0 ),
    .i1(\inst_dob_mux_b6/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b6/B0_2 ),
    .i1(\inst_dob_mux_b6/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b6/B0_20 ),
    .i1(\inst_dob_mux_b6/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_10 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b6/B0_22 ),
    .i1(\inst_dob_mux_b6/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_11 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b6/B0_24 ),
    .i1(\inst_dob_mux_b6/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_12 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b6/B0_26 ),
    .i1(\inst_dob_mux_b6/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_13 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b6/B0_28 ),
    .i1(\inst_dob_mux_b6/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_14 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b6/B0_30 ),
    .i1(\inst_dob_mux_b6/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_15 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b6/B0_32 ),
    .i1(\inst_dob_mux_b6/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_16 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b6/B0_34 ),
    .i1(\inst_dob_mux_b6/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_17 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b6/B0_36 ),
    .i1(\inst_dob_mux_b6/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_18 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b6/B0_38 ),
    .i1(\inst_dob_mux_b6/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_19 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b6/B0_4 ),
    .i1(\inst_dob_mux_b6/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b6/B0_40 ),
    .i1(\inst_dob_mux_b6/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_20 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b6/B0_42 ),
    .i1(\inst_dob_mux_b6/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_21 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b6/B0_44 ),
    .i1(\inst_dob_mux_b6/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_22 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b6/B0_46 ),
    .i1(\inst_dob_mux_b6/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_23 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b6/B0_48 ),
    .i1(\inst_dob_mux_b6/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_24 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b6/B0_50 ),
    .i1(\inst_dob_mux_b6/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_25 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b6/B0_52 ),
    .i1(\inst_dob_mux_b6/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_26 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b6/B0_54 ),
    .i1(\inst_dob_mux_b6/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_27 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b6/B0_56 ),
    .i1(\inst_dob_mux_b6/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_28 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b6/B0_58 ),
    .i1(\inst_dob_mux_b6/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_29 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b6/B0_6 ),
    .i1(\inst_dob_mux_b6/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b6/B0_60 ),
    .i1(\inst_dob_mux_b6/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_30 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b6/B0_62 ),
    .i1(\inst_dob_mux_b6/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_31 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b6/B0_8 ),
    .i1(\inst_dob_mux_b6/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_4 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b6/B0_10 ),
    .i1(\inst_dob_mux_b6/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_5 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b6/B0_12 ),
    .i1(\inst_dob_mux_b6/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_6 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b6/B0_14 ),
    .i1(\inst_dob_mux_b6/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_7 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b6/B0_16 ),
    .i1(\inst_dob_mux_b6/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_8 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b6/B0_18 ),
    .i1(\inst_dob_mux_b6/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_9 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b6/B1_0 ),
    .i1(\inst_dob_mux_b6/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b6/B1_2 ),
    .i1(\inst_dob_mux_b6/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b6/B1_20 ),
    .i1(\inst_dob_mux_b6/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_10 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b6/B1_22 ),
    .i1(\inst_dob_mux_b6/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_11 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b6/B1_24 ),
    .i1(\inst_dob_mux_b6/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_12 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b6/B1_26 ),
    .i1(\inst_dob_mux_b6/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_13 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b6/B1_28 ),
    .i1(\inst_dob_mux_b6/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_14 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b6/B1_30 ),
    .i1(\inst_dob_mux_b6/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_15 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b6/B1_4 ),
    .i1(\inst_dob_mux_b6/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b6/B1_6 ),
    .i1(\inst_dob_mux_b6/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b6/B1_8 ),
    .i1(\inst_dob_mux_b6/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_4 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b6/B1_10 ),
    .i1(\inst_dob_mux_b6/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_5 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b6/B1_12 ),
    .i1(\inst_dob_mux_b6/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_6 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b6/B1_14 ),
    .i1(\inst_dob_mux_b6/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_7 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b6/B1_16 ),
    .i1(\inst_dob_mux_b6/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_8 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b6/B1_18 ),
    .i1(\inst_dob_mux_b6/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_9 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b6/B2_0 ),
    .i1(\inst_dob_mux_b6/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b6/B3_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b6/B2_2 ),
    .i1(\inst_dob_mux_b6/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b6/B3_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b6/B2_4 ),
    .i1(\inst_dob_mux_b6/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b6/B3_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b6/B2_6 ),
    .i1(\inst_dob_mux_b6/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b6/B3_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b6/B2_8 ),
    .i1(\inst_dob_mux_b6/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b6/B3_4 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b6/B2_10 ),
    .i1(\inst_dob_mux_b6/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b6/B3_5 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b6/B2_12 ),
    .i1(\inst_dob_mux_b6/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b6/B3_6 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b6/B2_14 ),
    .i1(\inst_dob_mux_b6/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b6/B3_7 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b6/B3_0 ),
    .i1(\inst_dob_mux_b6/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b6/B4_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b6/B3_2 ),
    .i1(\inst_dob_mux_b6/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b6/B4_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b6/B3_4 ),
    .i1(\inst_dob_mux_b6/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b6/B4_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b6/B3_6 ),
    .i1(\inst_dob_mux_b6/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b6/B4_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b6/B4_0 ),
    .i1(\inst_dob_mux_b6/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b6/B5_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b6/B4_2 ),
    .i1(\inst_dob_mux_b6/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b6/B5_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b6/B5_0 ),
    .i1(\inst_dob_mux_b6/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[6]));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_0  (
    .i0(inst_dob_i0_007),
    .i1(inst_dob_i0_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_1  (
    .i0(inst_dob_i2_007),
    .i1(inst_dob_i2_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_10  (
    .i0(inst_dob_i20_007),
    .i1(inst_dob_i20_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_10 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_11  (
    .i0(inst_dob_i22_007),
    .i1(inst_dob_i22_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_11 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_12  (
    .i0(inst_dob_i24_007),
    .i1(inst_dob_i24_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_12 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_13  (
    .i0(inst_dob_i26_007),
    .i1(inst_dob_i26_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_13 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_14  (
    .i0(inst_dob_i28_007),
    .i1(inst_dob_i28_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_14 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_15  (
    .i0(inst_dob_i30_007),
    .i1(inst_dob_i30_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_15 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_16  (
    .i0(inst_dob_i32_007),
    .i1(inst_dob_i32_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_16 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_17  (
    .i0(inst_dob_i34_007),
    .i1(inst_dob_i34_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_17 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_18  (
    .i0(inst_dob_i36_007),
    .i1(inst_dob_i36_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_18 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_19  (
    .i0(inst_dob_i38_007),
    .i1(inst_dob_i38_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_19 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_2  (
    .i0(inst_dob_i4_007),
    .i1(inst_dob_i4_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_20  (
    .i0(inst_dob_i40_007),
    .i1(inst_dob_i40_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_20 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_21  (
    .i0(inst_dob_i42_007),
    .i1(inst_dob_i42_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_21 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_22  (
    .i0(inst_dob_i44_007),
    .i1(inst_dob_i44_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_22 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_23  (
    .i0(inst_dob_i46_007),
    .i1(inst_dob_i46_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_23 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_24  (
    .i0(inst_dob_i48_007),
    .i1(inst_dob_i48_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_24 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_25  (
    .i0(inst_dob_i50_007),
    .i1(inst_dob_i50_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_25 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_26  (
    .i0(inst_dob_i52_007),
    .i1(inst_dob_i52_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_26 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_27  (
    .i0(inst_dob_i54_007),
    .i1(inst_dob_i54_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_27 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_28  (
    .i0(inst_dob_i56_007),
    .i1(inst_dob_i56_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_28 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_29  (
    .i0(inst_dob_i58_007),
    .i1(inst_dob_i58_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_29 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_3  (
    .i0(inst_dob_i6_007),
    .i1(inst_dob_i6_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_30  (
    .i0(inst_dob_i60_007),
    .i1(inst_dob_i60_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_30 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_31  (
    .i0(inst_dob_i62_007),
    .i1(inst_dob_i62_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_31 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_32  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_32 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_33  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_33 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_34  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_34 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_35  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_35 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_36  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_36 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_37  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_37 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_38  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_38 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_39  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_39 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_4  (
    .i0(inst_dob_i8_007),
    .i1(inst_dob_i8_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_4 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_40  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_40 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_41  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_41 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_42  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_42 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_43  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_43 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_44  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_44 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_45  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_45 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_46  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_46 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_47  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_47 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_48  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_48 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_49  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_49 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_5  (
    .i0(inst_dob_i10_007),
    .i1(inst_dob_i10_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_5 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_50  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_50 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_51  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_51 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_52  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_52 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_53  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_53 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_54  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_54 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_55  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_55 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_56  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_56 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_57  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_57 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_58  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_58 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_59  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_59 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_6  (
    .i0(inst_dob_i12_007),
    .i1(inst_dob_i12_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_6 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_60  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_60 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_61  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_61 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_62  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_62 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_63  (
    .i0(inst_dob_i64_007),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_63 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_7  (
    .i0(inst_dob_i14_007),
    .i1(inst_dob_i14_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_7 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_8  (
    .i0(inst_dob_i16_007),
    .i1(inst_dob_i16_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_8 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_9  (
    .i0(inst_dob_i18_007),
    .i1(inst_dob_i18_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_9 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b7/B0_0 ),
    .i1(\inst_dob_mux_b7/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b7/B0_2 ),
    .i1(\inst_dob_mux_b7/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b7/B0_20 ),
    .i1(\inst_dob_mux_b7/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_10 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b7/B0_22 ),
    .i1(\inst_dob_mux_b7/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_11 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b7/B0_24 ),
    .i1(\inst_dob_mux_b7/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_12 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b7/B0_26 ),
    .i1(\inst_dob_mux_b7/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_13 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b7/B0_28 ),
    .i1(\inst_dob_mux_b7/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_14 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b7/B0_30 ),
    .i1(\inst_dob_mux_b7/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_15 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b7/B0_32 ),
    .i1(\inst_dob_mux_b7/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_16 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b7/B0_34 ),
    .i1(\inst_dob_mux_b7/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_17 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b7/B0_36 ),
    .i1(\inst_dob_mux_b7/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_18 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b7/B0_38 ),
    .i1(\inst_dob_mux_b7/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_19 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b7/B0_4 ),
    .i1(\inst_dob_mux_b7/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b7/B0_40 ),
    .i1(\inst_dob_mux_b7/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_20 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b7/B0_42 ),
    .i1(\inst_dob_mux_b7/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_21 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b7/B0_44 ),
    .i1(\inst_dob_mux_b7/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_22 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b7/B0_46 ),
    .i1(\inst_dob_mux_b7/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_23 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b7/B0_48 ),
    .i1(\inst_dob_mux_b7/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_24 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b7/B0_50 ),
    .i1(\inst_dob_mux_b7/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_25 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b7/B0_52 ),
    .i1(\inst_dob_mux_b7/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_26 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b7/B0_54 ),
    .i1(\inst_dob_mux_b7/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_27 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b7/B0_56 ),
    .i1(\inst_dob_mux_b7/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_28 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b7/B0_58 ),
    .i1(\inst_dob_mux_b7/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_29 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b7/B0_6 ),
    .i1(\inst_dob_mux_b7/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b7/B0_60 ),
    .i1(\inst_dob_mux_b7/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_30 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b7/B0_62 ),
    .i1(\inst_dob_mux_b7/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_31 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b7/B0_8 ),
    .i1(\inst_dob_mux_b7/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_4 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b7/B0_10 ),
    .i1(\inst_dob_mux_b7/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_5 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b7/B0_12 ),
    .i1(\inst_dob_mux_b7/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_6 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b7/B0_14 ),
    .i1(\inst_dob_mux_b7/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_7 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b7/B0_16 ),
    .i1(\inst_dob_mux_b7/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_8 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b7/B0_18 ),
    .i1(\inst_dob_mux_b7/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_9 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b7/B1_0 ),
    .i1(\inst_dob_mux_b7/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b7/B1_2 ),
    .i1(\inst_dob_mux_b7/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b7/B1_20 ),
    .i1(\inst_dob_mux_b7/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_10 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b7/B1_22 ),
    .i1(\inst_dob_mux_b7/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_11 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b7/B1_24 ),
    .i1(\inst_dob_mux_b7/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_12 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b7/B1_26 ),
    .i1(\inst_dob_mux_b7/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_13 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b7/B1_28 ),
    .i1(\inst_dob_mux_b7/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_14 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b7/B1_30 ),
    .i1(\inst_dob_mux_b7/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_15 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b7/B1_4 ),
    .i1(\inst_dob_mux_b7/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b7/B1_6 ),
    .i1(\inst_dob_mux_b7/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b7/B1_8 ),
    .i1(\inst_dob_mux_b7/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_4 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b7/B1_10 ),
    .i1(\inst_dob_mux_b7/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_5 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b7/B1_12 ),
    .i1(\inst_dob_mux_b7/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_6 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b7/B1_14 ),
    .i1(\inst_dob_mux_b7/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_7 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b7/B1_16 ),
    .i1(\inst_dob_mux_b7/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_8 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b7/B1_18 ),
    .i1(\inst_dob_mux_b7/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_9 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b7/B2_0 ),
    .i1(\inst_dob_mux_b7/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b7/B3_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b7/B2_2 ),
    .i1(\inst_dob_mux_b7/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b7/B3_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b7/B2_4 ),
    .i1(\inst_dob_mux_b7/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b7/B3_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b7/B2_6 ),
    .i1(\inst_dob_mux_b7/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b7/B3_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b7/B2_8 ),
    .i1(\inst_dob_mux_b7/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b7/B3_4 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b7/B2_10 ),
    .i1(\inst_dob_mux_b7/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b7/B3_5 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b7/B2_12 ),
    .i1(\inst_dob_mux_b7/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b7/B3_6 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b7/B2_14 ),
    .i1(\inst_dob_mux_b7/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b7/B3_7 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b7/B3_0 ),
    .i1(\inst_dob_mux_b7/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b7/B4_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b7/B3_2 ),
    .i1(\inst_dob_mux_b7/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b7/B4_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b7/B3_4 ),
    .i1(\inst_dob_mux_b7/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b7/B4_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b7/B3_6 ),
    .i1(\inst_dob_mux_b7/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b7/B4_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b7/B4_0 ),
    .i1(\inst_dob_mux_b7/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b7/B5_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b7/B4_2 ),
    .i1(\inst_dob_mux_b7/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b7/B5_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b7/B5_0 ),
    .i1(\inst_dob_mux_b7/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[7]));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_0  (
    .i0(inst_dob_i0_008),
    .i1(inst_dob_i0_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_1  (
    .i0(inst_dob_i2_008),
    .i1(inst_dob_i2_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_10  (
    .i0(inst_dob_i20_008),
    .i1(inst_dob_i20_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_10 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_11  (
    .i0(inst_dob_i22_008),
    .i1(inst_dob_i22_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_11 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_12  (
    .i0(inst_dob_i24_008),
    .i1(inst_dob_i24_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_12 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_13  (
    .i0(inst_dob_i26_008),
    .i1(inst_dob_i26_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_13 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_14  (
    .i0(inst_dob_i28_008),
    .i1(inst_dob_i28_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_14 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_15  (
    .i0(inst_dob_i30_008),
    .i1(inst_dob_i30_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_15 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_16  (
    .i0(inst_dob_i32_008),
    .i1(inst_dob_i32_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_16 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_17  (
    .i0(inst_dob_i34_008),
    .i1(inst_dob_i34_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_17 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_18  (
    .i0(inst_dob_i36_008),
    .i1(inst_dob_i36_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_18 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_19  (
    .i0(inst_dob_i38_008),
    .i1(inst_dob_i38_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_19 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_2  (
    .i0(inst_dob_i4_008),
    .i1(inst_dob_i4_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_20  (
    .i0(inst_dob_i40_008),
    .i1(inst_dob_i40_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_20 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_21  (
    .i0(inst_dob_i42_008),
    .i1(inst_dob_i42_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_21 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_22  (
    .i0(inst_dob_i44_008),
    .i1(inst_dob_i44_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_22 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_23  (
    .i0(inst_dob_i46_008),
    .i1(inst_dob_i46_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_23 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_24  (
    .i0(inst_dob_i48_008),
    .i1(inst_dob_i48_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_24 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_25  (
    .i0(inst_dob_i50_008),
    .i1(inst_dob_i50_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_25 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_26  (
    .i0(inst_dob_i52_008),
    .i1(inst_dob_i52_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_26 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_27  (
    .i0(inst_dob_i54_008),
    .i1(inst_dob_i54_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_27 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_28  (
    .i0(inst_dob_i56_008),
    .i1(inst_dob_i56_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_28 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_29  (
    .i0(inst_dob_i58_008),
    .i1(inst_dob_i58_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_29 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_3  (
    .i0(inst_dob_i6_008),
    .i1(inst_dob_i6_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_30  (
    .i0(inst_dob_i60_008),
    .i1(inst_dob_i60_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_30 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_31  (
    .i0(inst_dob_i62_008),
    .i1(inst_dob_i62_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_31 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_32  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_32 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_33  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_33 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_34  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_34 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_35  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_35 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_36  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_36 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_37  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_37 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_38  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_38 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_39  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_39 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_4  (
    .i0(inst_dob_i8_008),
    .i1(inst_dob_i8_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_4 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_40  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_40 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_41  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_41 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_42  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_42 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_43  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_43 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_44  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_44 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_45  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_45 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_46  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_46 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_47  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_47 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_48  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_48 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_49  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_49 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_5  (
    .i0(inst_dob_i10_008),
    .i1(inst_dob_i10_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_5 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_50  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_50 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_51  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_51 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_52  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_52 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_53  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_53 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_54  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_54 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_55  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_55 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_56  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_56 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_57  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_57 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_58  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_58 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_59  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_59 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_6  (
    .i0(inst_dob_i12_008),
    .i1(inst_dob_i12_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_6 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_60  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_60 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_61  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_61 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_62  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_62 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_63  (
    .i0(inst_dob_i64_008),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_63 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_7  (
    .i0(inst_dob_i14_008),
    .i1(inst_dob_i14_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_7 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_8  (
    .i0(inst_dob_i16_008),
    .i1(inst_dob_i16_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_8 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_9  (
    .i0(inst_dob_i18_008),
    .i1(inst_dob_i18_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_9 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b8/B0_0 ),
    .i1(\inst_dob_mux_b8/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b8/B0_2 ),
    .i1(\inst_dob_mux_b8/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b8/B0_20 ),
    .i1(\inst_dob_mux_b8/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_10 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b8/B0_22 ),
    .i1(\inst_dob_mux_b8/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_11 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b8/B0_24 ),
    .i1(\inst_dob_mux_b8/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_12 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b8/B0_26 ),
    .i1(\inst_dob_mux_b8/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_13 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b8/B0_28 ),
    .i1(\inst_dob_mux_b8/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_14 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b8/B0_30 ),
    .i1(\inst_dob_mux_b8/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_15 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b8/B0_32 ),
    .i1(\inst_dob_mux_b8/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_16 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b8/B0_34 ),
    .i1(\inst_dob_mux_b8/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_17 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b8/B0_36 ),
    .i1(\inst_dob_mux_b8/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_18 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b8/B0_38 ),
    .i1(\inst_dob_mux_b8/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_19 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b8/B0_4 ),
    .i1(\inst_dob_mux_b8/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b8/B0_40 ),
    .i1(\inst_dob_mux_b8/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_20 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b8/B0_42 ),
    .i1(\inst_dob_mux_b8/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_21 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b8/B0_44 ),
    .i1(\inst_dob_mux_b8/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_22 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b8/B0_46 ),
    .i1(\inst_dob_mux_b8/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_23 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b8/B0_48 ),
    .i1(\inst_dob_mux_b8/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_24 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b8/B0_50 ),
    .i1(\inst_dob_mux_b8/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_25 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b8/B0_52 ),
    .i1(\inst_dob_mux_b8/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_26 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b8/B0_54 ),
    .i1(\inst_dob_mux_b8/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_27 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b8/B0_56 ),
    .i1(\inst_dob_mux_b8/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_28 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b8/B0_58 ),
    .i1(\inst_dob_mux_b8/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_29 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b8/B0_6 ),
    .i1(\inst_dob_mux_b8/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b8/B0_60 ),
    .i1(\inst_dob_mux_b8/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_30 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b8/B0_62 ),
    .i1(\inst_dob_mux_b8/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_31 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b8/B0_8 ),
    .i1(\inst_dob_mux_b8/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_4 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b8/B0_10 ),
    .i1(\inst_dob_mux_b8/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_5 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b8/B0_12 ),
    .i1(\inst_dob_mux_b8/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_6 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b8/B0_14 ),
    .i1(\inst_dob_mux_b8/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_7 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b8/B0_16 ),
    .i1(\inst_dob_mux_b8/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_8 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b8/B0_18 ),
    .i1(\inst_dob_mux_b8/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_9 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b8/B1_0 ),
    .i1(\inst_dob_mux_b8/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b8/B1_2 ),
    .i1(\inst_dob_mux_b8/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b8/B1_20 ),
    .i1(\inst_dob_mux_b8/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_10 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b8/B1_22 ),
    .i1(\inst_dob_mux_b8/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_11 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b8/B1_24 ),
    .i1(\inst_dob_mux_b8/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_12 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b8/B1_26 ),
    .i1(\inst_dob_mux_b8/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_13 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b8/B1_28 ),
    .i1(\inst_dob_mux_b8/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_14 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b8/B1_30 ),
    .i1(\inst_dob_mux_b8/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_15 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b8/B1_4 ),
    .i1(\inst_dob_mux_b8/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b8/B1_6 ),
    .i1(\inst_dob_mux_b8/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b8/B1_8 ),
    .i1(\inst_dob_mux_b8/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_4 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b8/B1_10 ),
    .i1(\inst_dob_mux_b8/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_5 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b8/B1_12 ),
    .i1(\inst_dob_mux_b8/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_6 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b8/B1_14 ),
    .i1(\inst_dob_mux_b8/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_7 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b8/B1_16 ),
    .i1(\inst_dob_mux_b8/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_8 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b8/B1_18 ),
    .i1(\inst_dob_mux_b8/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_9 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b8/B2_0 ),
    .i1(\inst_dob_mux_b8/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b8/B3_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b8/B2_2 ),
    .i1(\inst_dob_mux_b8/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b8/B3_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b8/B2_4 ),
    .i1(\inst_dob_mux_b8/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b8/B3_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b8/B2_6 ),
    .i1(\inst_dob_mux_b8/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b8/B3_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b8/B2_8 ),
    .i1(\inst_dob_mux_b8/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b8/B3_4 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b8/B2_10 ),
    .i1(\inst_dob_mux_b8/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b8/B3_5 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b8/B2_12 ),
    .i1(\inst_dob_mux_b8/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b8/B3_6 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b8/B2_14 ),
    .i1(\inst_dob_mux_b8/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b8/B3_7 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b8/B3_0 ),
    .i1(\inst_dob_mux_b8/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b8/B4_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b8/B3_2 ),
    .i1(\inst_dob_mux_b8/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b8/B4_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b8/B3_4 ),
    .i1(\inst_dob_mux_b8/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b8/B4_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b8/B3_6 ),
    .i1(\inst_dob_mux_b8/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b8/B4_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b8/B4_0 ),
    .i1(\inst_dob_mux_b8/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b8/B5_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b8/B4_2 ),
    .i1(\inst_dob_mux_b8/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b8/B5_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b8/B5_0 ),
    .i1(\inst_dob_mux_b8/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[8]));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_0  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_1  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_10  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_10 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_11  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_11 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_12  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_12 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_13  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_13 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_14  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_14 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_15  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_15 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_16  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_16 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_17  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_17 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_18  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_18 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_19  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_19 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_2  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_2 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_20  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_20 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_21  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_21 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_22  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_22 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_23  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i32_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_23 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_24  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_24 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_25  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_25 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_26  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_26 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_27  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_27 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_28  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_28 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_29  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_29 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_3  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_3 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_30  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_30 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_31  (
    .i0(inst_dob_i48_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_31 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_32  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_32 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_33  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_33 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_34  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_34 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_35  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_35 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_36  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_36 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_37  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_37 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_38  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_38 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_39  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_39 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_4  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_4 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_40  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_40 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_41  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_41 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_42  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_42 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_43  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_43 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_44  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_44 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_45  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_45 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_46  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_46 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_47  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_47 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_48  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_48 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_49  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_49 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_5  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_5 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_50  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_50 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_51  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_51 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_52  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_52 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_53  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_53 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_54  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_54 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_55  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_55 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_56  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_56 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_57  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_57 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_58  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_58 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_59  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_59 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_6  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_6 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_60  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_60 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_61  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_61 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_62  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_62 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_63  (
    .i0(inst_dob_i64_009),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_63 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_7  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i0_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_7 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_8  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_8 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_9  (
    .i0(inst_dob_i16_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_9 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b9/B0_0 ),
    .i1(\inst_dob_mux_b9/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b9/B0_2 ),
    .i1(\inst_dob_mux_b9/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_10  (
    .i0(\inst_dob_mux_b9/B0_20 ),
    .i1(\inst_dob_mux_b9/B0_21 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_10 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_11  (
    .i0(\inst_dob_mux_b9/B0_22 ),
    .i1(\inst_dob_mux_b9/B0_23 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_11 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_12  (
    .i0(\inst_dob_mux_b9/B0_24 ),
    .i1(\inst_dob_mux_b9/B0_25 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_12 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_13  (
    .i0(\inst_dob_mux_b9/B0_26 ),
    .i1(\inst_dob_mux_b9/B0_27 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_13 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_14  (
    .i0(\inst_dob_mux_b9/B0_28 ),
    .i1(\inst_dob_mux_b9/B0_29 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_14 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_15  (
    .i0(\inst_dob_mux_b9/B0_30 ),
    .i1(\inst_dob_mux_b9/B0_31 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_15 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_16  (
    .i0(\inst_dob_mux_b9/B0_32 ),
    .i1(\inst_dob_mux_b9/B0_33 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_16 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_17  (
    .i0(\inst_dob_mux_b9/B0_34 ),
    .i1(\inst_dob_mux_b9/B0_35 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_17 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_18  (
    .i0(\inst_dob_mux_b9/B0_36 ),
    .i1(\inst_dob_mux_b9/B0_37 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_18 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_19  (
    .i0(\inst_dob_mux_b9/B0_38 ),
    .i1(\inst_dob_mux_b9/B0_39 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_19 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_2  (
    .i0(\inst_dob_mux_b9/B0_4 ),
    .i1(\inst_dob_mux_b9/B0_5 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_2 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_20  (
    .i0(\inst_dob_mux_b9/B0_40 ),
    .i1(\inst_dob_mux_b9/B0_41 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_20 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_21  (
    .i0(\inst_dob_mux_b9/B0_42 ),
    .i1(\inst_dob_mux_b9/B0_43 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_21 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_22  (
    .i0(\inst_dob_mux_b9/B0_44 ),
    .i1(\inst_dob_mux_b9/B0_45 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_22 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_23  (
    .i0(\inst_dob_mux_b9/B0_46 ),
    .i1(\inst_dob_mux_b9/B0_47 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_23 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_24  (
    .i0(\inst_dob_mux_b9/B0_48 ),
    .i1(\inst_dob_mux_b9/B0_49 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_24 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_25  (
    .i0(\inst_dob_mux_b9/B0_50 ),
    .i1(\inst_dob_mux_b9/B0_51 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_25 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_26  (
    .i0(\inst_dob_mux_b9/B0_52 ),
    .i1(\inst_dob_mux_b9/B0_53 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_26 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_27  (
    .i0(\inst_dob_mux_b9/B0_54 ),
    .i1(\inst_dob_mux_b9/B0_55 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_27 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_28  (
    .i0(\inst_dob_mux_b9/B0_56 ),
    .i1(\inst_dob_mux_b9/B0_57 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_28 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_29  (
    .i0(\inst_dob_mux_b9/B0_58 ),
    .i1(\inst_dob_mux_b9/B0_59 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_29 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_3  (
    .i0(\inst_dob_mux_b9/B0_6 ),
    .i1(\inst_dob_mux_b9/B0_7 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_3 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_30  (
    .i0(\inst_dob_mux_b9/B0_60 ),
    .i1(\inst_dob_mux_b9/B0_61 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_30 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_31  (
    .i0(\inst_dob_mux_b9/B0_62 ),
    .i1(\inst_dob_mux_b9/B0_63 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_31 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_4  (
    .i0(\inst_dob_mux_b9/B0_8 ),
    .i1(\inst_dob_mux_b9/B0_9 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_4 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_5  (
    .i0(\inst_dob_mux_b9/B0_10 ),
    .i1(\inst_dob_mux_b9/B0_11 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_5 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_6  (
    .i0(\inst_dob_mux_b9/B0_12 ),
    .i1(\inst_dob_mux_b9/B0_13 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_6 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_7  (
    .i0(\inst_dob_mux_b9/B0_14 ),
    .i1(\inst_dob_mux_b9/B0_15 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_7 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_8  (
    .i0(\inst_dob_mux_b9/B0_16 ),
    .i1(\inst_dob_mux_b9/B0_17 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_8 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_9  (
    .i0(\inst_dob_mux_b9/B0_18 ),
    .i1(\inst_dob_mux_b9/B0_19 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_9 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b9/B1_0 ),
    .i1(\inst_dob_mux_b9/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b9/B1_2 ),
    .i1(\inst_dob_mux_b9/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_10  (
    .i0(\inst_dob_mux_b9/B1_20 ),
    .i1(\inst_dob_mux_b9/B1_21 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_10 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_11  (
    .i0(\inst_dob_mux_b9/B1_22 ),
    .i1(\inst_dob_mux_b9/B1_23 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_11 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_12  (
    .i0(\inst_dob_mux_b9/B1_24 ),
    .i1(\inst_dob_mux_b9/B1_25 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_12 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_13  (
    .i0(\inst_dob_mux_b9/B1_26 ),
    .i1(\inst_dob_mux_b9/B1_27 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_13 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_14  (
    .i0(\inst_dob_mux_b9/B1_28 ),
    .i1(\inst_dob_mux_b9/B1_29 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_14 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_15  (
    .i0(\inst_dob_mux_b9/B1_30 ),
    .i1(\inst_dob_mux_b9/B1_31 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_15 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b9/B1_4 ),
    .i1(\inst_dob_mux_b9/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_2 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b9/B1_6 ),
    .i1(\inst_dob_mux_b9/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_3 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b9/B1_8 ),
    .i1(\inst_dob_mux_b9/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_4 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b9/B1_10 ),
    .i1(\inst_dob_mux_b9/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_5 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b9/B1_12 ),
    .i1(\inst_dob_mux_b9/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_6 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b9/B1_14 ),
    .i1(\inst_dob_mux_b9/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_7 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_8  (
    .i0(\inst_dob_mux_b9/B1_16 ),
    .i1(\inst_dob_mux_b9/B1_17 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_8 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_9  (
    .i0(\inst_dob_mux_b9/B1_18 ),
    .i1(\inst_dob_mux_b9/B1_19 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b9/B2_9 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b9/B2_0 ),
    .i1(\inst_dob_mux_b9/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b9/B3_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b9/B2_2 ),
    .i1(\inst_dob_mux_b9/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b9/B3_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b9/B2_4 ),
    .i1(\inst_dob_mux_b9/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b9/B3_2 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b9/B2_6 ),
    .i1(\inst_dob_mux_b9/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b9/B3_3 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_4  (
    .i0(\inst_dob_mux_b9/B2_8 ),
    .i1(\inst_dob_mux_b9/B2_9 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b9/B3_4 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_5  (
    .i0(\inst_dob_mux_b9/B2_10 ),
    .i1(\inst_dob_mux_b9/B2_11 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b9/B3_5 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_6  (
    .i0(\inst_dob_mux_b9/B2_12 ),
    .i1(\inst_dob_mux_b9/B2_13 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b9/B3_6 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_3_7  (
    .i0(\inst_dob_mux_b9/B2_14 ),
    .i1(\inst_dob_mux_b9/B2_15 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b9/B3_7 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b9/B3_0 ),
    .i1(\inst_dob_mux_b9/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b9/B4_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b9/B3_2 ),
    .i1(\inst_dob_mux_b9/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b9/B4_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_4_2  (
    .i0(\inst_dob_mux_b9/B3_4 ),
    .i1(\inst_dob_mux_b9/B3_5 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b9/B4_2 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_4_3  (
    .i0(\inst_dob_mux_b9/B3_6 ),
    .i1(\inst_dob_mux_b9/B3_7 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b9/B4_3 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b9/B4_0 ),
    .i1(\inst_dob_mux_b9/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b9/B5_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_5_1  (
    .i0(\inst_dob_mux_b9/B4_2 ),
    .i1(\inst_dob_mux_b9/B4_3 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b9/B5_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b9/B5_0 ),
    .i1(\inst_dob_mux_b9/B5_1 ),
    .sel(addrb_piped[6]),
    .o(dob[9]));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

