module sync( );



endmodule
